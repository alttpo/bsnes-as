BSV1n BST1108.4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �7�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    � �                                                                                                                                                                                                                                                                                                                                                                       �                                                                                                � � � � � �U                              ��                                                                                                                                                                                                                                                       �l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ i�    ��  �            ��   ~ B~   ��G            T  �   ,     T  l5    t k6        �  5 l�� � �               5l ��           x      	                     ��             0        d9
	    � @�             $  ��
  �  ~ ~ ~�� 2� ~� ~� ~ !~�!~ "~          �                0�     B       ^                        ;                                                                                                                     �  "� ����������������   � ��� ����P ���ʨȵ���@�       �26�     '     �      � K @`  AH ��                                                                                                                                                               @ 	       �    @     $`  p0                                                                                                          �
                           �                    P         H{    �	               �                                                                                               0�                     ��                                      0 +    p                              T# p              %                �                                                                                                  � � � �                         P&P(,(,*                        �                  �                  MMMMMM�                  MMMMMM�                       x          P   @                       x z �     ����                                                                   �   E 3    ~               �              �               �    �	�2  �;            �               ���      �
                  6        �� ~       �           � @                                                                                                                                                                                                                        ��`8��88x�88�� ��� ��� =�� }�� ��� ���4;0�=8�=��4��4��88��$���m���mh������-m𛤀��= ��=���=P`�= P�=G�[�dG�$J�-]��e�$b�dZ�'��l���"���"���"v�l���"}��"x��"s��"w�lq�lq�ln�l��Fv� (v�"hK�[�k�{�K��[����n0�.v� .v�.��*�� n��n{�*(�7=0�8=v�l(~�lh|� h|�"h8�8�@�7�(�7=0�8=8�8=@�7}(�7�0�8�8�8�@�7���D��D��g��f��}��m��~��n��nT�BYU�BYb�Yx� (x�"he� (e�"hr�&dI�MY<�l;�l��*���dk6 .l=.�� .j� .j�.t:*��.��*mFl(uFlhl4 hl>"hc� hc�"hx� x� ��,1��q��1��1x�l(��+�� )��+ �   �  �� ��
( ������
  � (�������
                                                F
          
           �����@���@� � �@�@�@�@�������  �� �    @ � ����@�@�  @�@�        ������� ������p                                                   �   ��              ha        ! "  0000000000(  00                    	                 �����������������?������������� ���  �         b  �� �  I8  ?�    #!       	          �             �   �        ��    �                     $                               0  00    0       !!�!                                                               >   P`���pp����P�@�C P� ��P� ���)�                                             � �             � @                          	                                                  									                                                                   mmmmmmm�m?K���                     ��  ���� ��   AA�]���                           �                                                                                                                                                                            �     MBL     CC  D  DD�                       �    ��         �     � z       P�� r     �����    l5                  P     h �  0  @                      <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�(�(���������H<<<<<<<<<<<<<<<<<<<<<�(�(��������H�H<<<<<<<<<<<<<<<<<<<<<�(�(�������H�H�H<<<<<<<<<<<<<<<<<<<<<-h,h�������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H���������H<<<<<<<<<<<<���������H�H���������H�H<<<<<<<<<<<<���������H���������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<�Ȱ�����������������H�H�H<<<<<<<<<<<<�����������������������������������șH�H<<<<<<<<<<<<�������������������������������������ȒH<<<<<<<<<<<<����������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�Y��Y�����������������5�5�5�5�5�5�5�u�ub �5�5d@4t �u�u� �5�5�@4� �u�u� '�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�u�u� '�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�u�u� �5�@2�5� �5�"�5�"�5B �5C@2�5] �5@24#@24C@24c@24�@24�@24�@24�@24@24#@24C@24c@24�@24�@24�@24�@24@24#@24�                                             D @              @	            �;�3              �+                                                                          5          l���������}}~~��xx                    		                                                                                                                                         � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                %a%a    Z  9P   �9          )                               mmoo�mmmm�m?K���dhs��������)�  ��Os<����P�@�C       	   	                     M�		M  BL    0    0(  00           ��  ���                         		��  ���       ��                     ` P     K_u Lo          �p�     X0X �|                                                                                                                                                                                        � 1                          /�/�~ & 
/�	     2�	 ���� (
   �   @   @       @  3 4                                  3344                                    �   
�      34                       �44���44� �             <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<���������������������������������������������H<<<<<<<<<<<<<<<<<<<��������������������������������������������H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<�������������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<������������������,�-�-�,����������������������H�H�H<<<<<<<<<<<<<<<<<<<�����������������������������������������������������������������������������������șH�H<<<<<<<<<<<<<<<<<<<��������������������������������������������������������������������������������������ȒH<<<<<<<<<<<<<<<<<<<������������������������������������������������������������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<����������(�(�(�(���������H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<����������(�(�(�(��������H�H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<����������(�(�(�(�������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<���������,(-(-h,h�������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<��������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<��������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�����������������������������H�H�H���������H<<<<<<<<<<<<<<<<<<<<<<<<�����������������������������H�H���������H�H<<<<<<<<<<<<<<<<<<<<<<<<�����������������������������H���������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<�����������������������Ȱ�����������������H�H�H<<<<<<<<<<<<<<<<<<<<<<<<�������������������������������������������������������������������������șH�H<<<<<<<<<<<<<<<<<<<<<<<<����������������������������������������������������������������������������ȒH<<<<<<<<<<<<<<<<<<<<<<<<��������������������������������������������������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������8�8�8�8�8��������������������������������FPQPPQPQPQPQPQPQPQPQPQPQPQPQ(P(Q(P(�(�(�h�hQ(PQFH�������������������������CGa``a`a`a`a`a`a`a`a`a`a`a`a(`(a(`((�	�	ha`GHCH�������������������������STHppppppppppppppppppppppppp(p(p(p((HpHHTHSH�������������������������CDq��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P�PqHDHCH�������������������������CDq�����������������������������������qHDHCH�������������������������STq����������������������((M���������PqHTHSH�������������������������CDq�����������������������88M����������qHDHCH�������������������������STq���������������������������������PqHTHSH�������������������������CDq�����������������������������������qHDHCH�������������������������STq����((M����������������((M���������PqHTHSH�������������������������CDq�����88M����������������88M����������qHDHCH�������������������������STq���������������������������������PqHTHSH�������������������������CDq�����������������������������������qHDHCH�������������������������STq����((M���������������������������PqHTHSH�������������������������CDq�����88M����������������������������qHDHCH�������������������������STq���������������������������������PqHTHSH�������������������������STq���Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ю�qHTHSH�������������������������CDH�p�p�p�p�p�p�p�p�p�p�p�p��x�x��p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�H�DHCH�������������������������SG�a�`�`�a�`�a�`�a�`�a�`�a�`���	�	�a�`�a�`�a�`�a�`�a�`�a�`�a�`�a�`�a�`�G�SH�������������������������F�P�Q�P�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�F��������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H����������������������������������������������������FPQPPQPQPQPQQPQFH������������������������������������������������CGa``a�	�	H`aa`GHCH������������������������������������������������STHpppxxHHpppHHTHSH������������������������������������������������CDq��P��P��P��P��PqHDHCH������������������������������������������������CDq������������qHDHCH������������������������������������������������STq����������PqHTHSH���������������������������������������FPQPPQPQPVTq����������PqHTHVHPQPQPQPQFH������������������������������CGa``a`a`aWq������������qHWH``a`a`a`GHCH������������������������������STHppppppppX����������PXHppppppppHHTHSH������������������������������CDq��P��P��P��P�����������P�P��P�P��P��P�PqHDHCH������������������������������CDq������������������������������qHDHCH������������������������������STq����������������������������PqHTHSH������������������������������CDq������������������������������qHDHCH������������������������������STq����������������������������PqHTHSH������������������������������CDq������������������������������qHDHCH������������������������������STq����������������������������PqHTHSH������������������������������STq���Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь���qHTHSH������������������������������CDH�p�p�p�p�p�p�p�p�p�p�p�p��5�5��p�p�p�p�p�p�p�p�p�p�p�p�H�DHCH������������������������������SG�a�`�`�a�`�a�`�a�`�a�`�a�`�$�%�%�$�a�`�a�`�a�`�a�`�a�`�a�a�`�G�SH������������������������������F�P�Q�P�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�Q�P�Q�F�������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������L�H�H�H��������������������������������������������������������������̥H�H�H�������������������������������������������������������������������������������������������� � � � � � � � �                                 � � � � � � � �         � � � � � � � �        ����������� �����   � � � � �����        � � � � � � � � ��������� � � �  7 M � ����������6�{rͺ�K���߷{����
�)� ���� � �������� �<�<� �=������<BB=�$!>�� � ��������Ab�                                                                                                �������������� ��������  � � � � � � � �                                                                                                                                                        �<�v�2�2�^�X�p�P�v22^YsW� �B��0���� ���;���� !�?�?�?�� � ��!@@@!> `d � sm^��ޛp���!!!                                                                                                                        �&� � �<� �~�~� XZBB~   � �`��?�?���  @@   �B�$�f�f�f�f�f�~ � 	w��ϼۼ[�[� ������[�I�d�0ϼ�����������ؿ�@������V�V�F�Z  QIIIE� � �?�0�!�,�$�0 @O^S[O����������       ?���                                                                         �  g{g � ������  � ��8���8��� � �      �8�\�m�~�}�{�&|�A!   8��<�x��D?Ŀa��8�                                                                                                                                                  �W�Z�_�o�w�8�� HE@`px � �&�6� ��U�?�@_YI  @??  � � � � � � ��������                                                                         � ��8���8��� � �       �  g{g � ������ ���?����?=���<   �  �`�k������Ө�Iv !"$@���B�N�f�:e�>�w�`1	 � �{�w�b�F�Q�Q�R D�|���}��|�9�����     O����������L�}��������  �� �m�j�m�v�j�j   ���0Oϰ�@���  0@�  � ��@�@�@�@�@�@ `````�  �  � � � � �  ��     �?��y��=�}�u��  
z?�_��s�y��l�l�d    p  ��?���_��?�? � ��x�s�g�o�o�o   ������������������������������������������������ ���|�{�w��     � � � � � � �� ���������M�!�A��6�6�U�A @*II*���k��x�i��2�V  `  �A�I�+�^�c�?�@�     @? �X_���?����     � �Y�Y�Y�Y�Y�Z�Z�T��3�'�/�/�/Я�        �@�@�@�@�@�@�_�@`ooooo� � � � � �  �   ����������������������
;????�`�`�f�f�F�c�8� / �_�_�O��?���o �c�`�p�x����      �^�F�w�u�z���     ��������������������������������         � ��g�N�]�{�w�n        � �o�i�i���� `f`````� �o�n�n���� `a`````� � � � � � � �  �  ����� ��������K�W�\�B�[�]�J�l Wh��Oϐp����p�@0���� �7�0�0�>�?�  00>>?  �� 	�	���  �� �  � � �{�t�d�D�S�P�X � �@�_�_�_�@��@ ?   ?                  ��������        �oP� ���W�k�k�c     ����������������        ���?��� � � �         �����������?��        ��	�o�i�o�v�I�O`f```pyO���o�n�o��`�`a```���� � � ����� xp`  ����������� ���  �g�s�y�|�~�7��      Hp ��5��������      �;�a�@��1�`�0� >`N����������    ���V�C�b�p�x���     �^�\�Y�S�G�@��       ? ?   � �         ���?�?������        �g�k�l�w�h�_��     � � � � � � � �         � ?                   � � � � � ?           ��������        ���6�����v�����        ��/������ � � ��    o��������������������8�����x�<���       `�l� � �w�������       ��������  ??��������  @???  ��������� ���C�y�|�~߿����;������������Ii�ͻ����F�  �(�W��� �@`�>�'o`? �#U�t�0Po��� �p���  À�x�~��b��� ?x�����@� � ��  �/��     ���� �� � �      j��� �� �� �     �� �����o�w�8�? @@�p�{�;� �  � � �p{;     ��������������������������r:���:_�U�U��*����8        �:�u�7���55  ��  �����@�?���`��_�??      � �������@�     N�����ֵŦäۼää���������[�kֹeھG���3    ���
6�� ;����p�  �2���6�,��51�2��'�������c � ���<>~�����*ށu+��Ww߯� �`����  ���/�[�3�}��p`@     �� �� 2��m�-� �   M   ��������   � � �������`�����e ����� � ���     77� � ��=�9�0� �   =90&/U��*�
?���|��       ����� ��� � ��� n`~� �?�?�?�?�?�?�? ?�� ������ ����Y ääääۼääѲ���������d����|� � �   ������  ��  �� ���       ���:���7�	  
�n�gjwvwrwr;9���������/h/hH��G�������00p`� ���~�A��~�A  <  <  ���<�{�~�}�{�w  �  ������  �����  ��  ��������������������������                                                ��K�x�{�x�x�0� x0      ��������       ��~�@���	��<      �o� ����� �m�m    @  ȹļ�������������������� `�?@������ ?��    � ������ �  �(((�  � ������ �  ����|}xy�y`a;��������� ��� ���� �  �   �� �`�`���� �p `ogsx�p���1���� ~~7;;;OH��_��	>?�  0����� �8�g������k� 8p  ��������pppppppp|������� ������|�w��w�w�w�7� � ������p?� � � � ����� � ??� � � � � � � � �������� �B���X��?����      � �P�i�>��/�w�v     �w�v�v�v�w�w�v�v   ������o�`�@��  O� � � � �    ��� ?��  �? ��E�U�Q�Y�M�E�U�Q:*.&2:*.� ��Q�Y�M�E�U�Q  .&2:*.m��?�O�o�q�~�w�w     � ߿��7�������{      �����އ�������� >><  �΋�OH��H��	��0p�0�p� � � �  � � � � ���    � � �    � � ��  ���    ��������pppppppp� � � � ����� �?� � � � � � � � ���������������������������������w�w�w�v�v�v�o�o     �o�o�k�m�W�'��    � ��hw�  ��� �   � �   �����P�V�D�E�Q�U?0/);:.*�T�V�@�F�@��� +)?9?     ss��  ����� ���1�   �!�s�y�|�|�?��        c� � ��   �� ��    �   �2��6M����� 0�   ��v��}�n��� �    �  ��������������������߿c�3��{vvvvv����� ���?p�?� ����   ���  ��������������������߿����7�o?��������߿������������������������                                                �x���p�� �@�~� x�p    �~�~�~�~�~�~�~�~        ����s缳߹o�w�wh�s��oww���<{Ͻ��{���s��<��{���                                                                                                                                                                                                                                                                                                                                                                                                �������������������߿�������������������߿�������������������߿�������������������߿�������������������߿�������������������߿                           � �       �          P l{4     p|w         
6�,    >�     337  ???    � ��~D;����  �4��g   
      � �`��,�p_�� ��vr���   > ?OKX  � ��0�<���� �� ������:�������������������߿�������������������߿�������������������߿�������������������߿�������������������߿�������������������߿        � ����x|8|8|   ����||| �c�h�	��n} �����=���� �l�r�|| �??���|7?   ?? � ����0p�� 0 �m"b���03?/& ??3:���l���`� �     ������  ��A�dw	> �z/���^ |0 � �}������   /7s ;,O  � ��0�8�����0 �����4�   ?7 #*  � `�x������8�p ������r          P l�t     p|�         
6�.    >�          0 H0w     0x         
�    �            8 '      8?           4�0     <�            8 '      8?           4�0     <� 0g8�p�`� �        � ��������     �8�?�8�;�;�;��    �4�����������    ���� ���`0? ��H6�y�����p��� �	l�0�3?77]8 -8/,z'� � � | ���p��� ����d�0��c�(�I�L}- ����?=��m��4�x�x�pp �??{���p�s�@�{7< ���O?<���<
�4����� �>������K5V)v	[$j4; GOo?��x�x��z\�0�� ��������M3Y'w7/	 GO;9� ���t��ĸ�0�� ���������9�
�e�b�a�p�8�8      ��y��C�`^�*ՙf�7       W/X'_ [$K4c0         ���������        <6>}"???~� ��� �0��(�8����x<l|> 8 ; lE:L7,(+__~?    � r̹n�.�v�  ��?� :~?� @��@� ��(�|�.؀����،�   /s,]n) 1]W~ �B�������~��~�~�������     /3}"  1=_  ~ �B�������~�� ~������    � ������0�D  ��Ȍ��      /3  1=  ~ �B�������~�� ~������       , < $ 4    4<<,        ` � ��    `���           ��(     �<^#! 7 {y>z������X0�� ��ޞ|�p�??_ 0w(: ??sO_?.�����,�p|���� ����|���_/.~=< ?���t~�<����0�@� ��������17    K; $����ý�<~�<�� �����~<�^o)?  gW+~�$�����=g��X� �������z�����@Ȱ� �   ������� =o-/';: /S3;'&~�$����ý�<�� �������444 $        ,,,<   ?_%L0~ ?  ?~s2<�������@� 0�� ��>~��0�        ` � ��    `���           ��(     �<        @ � ��     @���          p �0�P     p�x     ={$_O	  #]gw        ~ �~��<�    ~���       ={$_   #]g          ~ �~��     ~��      0 X �@�$�   0hĺ�8 < z4][O /	 <Nkm7      p �p�~?���   p���� 8  T T |                D � D                  < f$�B� �    <Z��� 8 llllll(TTTTTT    ?  �? ?     ?@�@? ?_%L0~ ?    ?~s2 <�������@��p� ��>~������~}3{A>> ���{A>x��h�X~������   ������� /	    7 �����<~��~�<<�� ������<�O	/	    w7 <������;{�ƽ�? �������?����@P��  �� � ����� ��           ���?�α�= �����8 (((((((8(((((((      � ��        ���  �$��Z $      ���f<  | T(D8(| D8( Dl|8|D(    � �d�6�d�     �z9z�      /?^#_1  77{     (�0��z���  8����       /   7       (�0��x�   8���   / 7   (�0��p����� 8���и / 7??    � ���������  ������     =6  ?    � � � ����m8  �����     =6  ?    � �`�0����}8  �����   //7 >?/      � p�8��(��   �����  ??~7?;w� ��� `���� �����������m�C��K     ����O
 ������u@� p     �����P  ?''36 ;=???�����̸l8�0x0 ܼ����x073   ?? ��̸�p�p�0p     �����p  ;7	 7?�0��x��������� ���ذ���'�o�~     w��  �<�|�������     ������  '�o�~       w��   �<�~���88       ����8   .?	?	?   ?;9- t������������   �؜���� |??     ? �x������ݸ�t`� ��������                                                  ??~7?;w� ��� `���� ����������  7';9  � � ��:�~��� �����ޜ .'/???� ��p�8�t����xx��������� ?2�c�g|?~?��    � � @�@�@��   ������ ?13>??ys??  � ���  � � �@� �������   <x��� 3W���  � ��|0�O   �0�
���      ` �`�`�@   `���       ���   ��                                                |??     ? �x�|�����8�t`� ��������/.   =?��t���� p@� � � ���а�`�7 ?x�p���8�p�� ��� ��������O~? _Ow'� ����m����   ������ ??'> /'?;� |8n<�t��5���� �|~������w5:;  �J/$�T �����  �Z�d�n=n;>8     ?8  v�v�<����       ��<��   �m�a�]�>����]eA>]���k��x�i��6�V��r`T�`�s�_�o�?e>	w,`3WO'	$    ? ??=;?   @ � x > =   	 @�X&#    � �0�:�y�� �����  c �  ?    ? � �f�B�f�<� � �  fJf���   ( ( h h h �   000p  4 : z z } �  <<>~  8?????? 8??????      ����������   �����                           ����      ��1111! !//   L L L L � ���xt8�����  ��I�I�+�^�c��� II*\@ �X_���?����� PB
��     ���  ���      � ��   ??� ?? {??G?����?�����o��y���������      ? � >       ?       � ~<= � �     ��� � � ����� � p`PPPP`p� ������� pnZPTZnp????1     ????1   �����������<� �����<            �����������     �����   /�_� �@      ? �8� � ~ ��� �� ������ �������������������߿<<B~�ý��[g~Z$$<~���gZ$�$�$�$�$�$�$�$�$ZZZZZZZZ,,vF����nn<< \8   204z   E� ��8 <0< ��  �����Bǂ�B@?@?�?����?�B" ��A�B��������ABDH ��� 8?8?????????� �����<����x�8��������                    ������     ���            ? �;���������� ?� �?�?�?�?��!^�� @H^!  �� � ���䅄{�  ��z� �������������������߿�$�$�$�$�<�~ < ZZZZBf< 8 D8�|��f~,<  8|f, 4,4,4,4,4,4,4,4,,,,,,,,,��Lo0 ~?  ��{~S/����� ~�� x�� ��~�������@?@?@?�_���� "B���������A�@�� DBA@?=???> ??????�8�x�x�x�xl���� ��������           �����������00   �����0  ???x8`  k6k6  @G_ww������
����@ @ @                                                                  000` `      > 7 3 a `          � � �           ���  <              <              � ��|88     ���D|(8    @ ` ` p 0 0      @ ` ` p 0 0     <(8        < 8 8   } � �           } � �                                 �               �                      0            0       � �� � � �      � � � � � �   < ~<<      $<B~$<   ` � � � � �   � ` � � � � �   �||�pp         |D|��pp                                       ��     ��  8   ?>      8!?">                      � � �`���       P��� ���    0             ?             ��|x00     ��D|Hx00     @   �           @   �          ` x |�X�pp      `x|����pp                                 �  ��          ������                             � 0 �           ������                             � @�@           ������


          P�P�P���@ �     ������������             ��� �@��     ������������                @ @ @�@��       ����������                           � � �0�� �     ��T�������� , f$~$� � ~ < 4<Z~Z~����~~$<$ ~ �n$f$�~ $ $$Z~��R~Z~��Z~$$     < < < < <     $<$<$<$<<<` � �� � �� ` ``������������``         $ ~$~$        <<Z~B~                 � �             H���            < < < < <      $<$<$<$<$<       , f$~$� � ~   4<Z~Z~����~~~ � ��$~$<     f~������B~<<        ?   ?         ??@@??    � � ~ < < <    ����f~$<$<$<                   � 0�h�8���    ��0�8����< B<�~�N�^�~�~B<<<Z~����������B~< B<B<R,B<B<B<< <<B~B~J~Z~B~B~<<   $< B<�~�<�B  <<<<B~������| �d�t�r�z�t�|| ||������������||      < B<�~�<�@      <<B~������             �``           ���``          $$$$$     <<<<<<<<<<     f�f�D�^�~�~~ ~~����������~~�~�f�f�~B<<     ��������B~<<                      �~�~�B�Zf$$ ��������~~<<<<                               ((T�(  (88\�(8 .R R �@�@�@,>PrPr����  1 N11       !1N1?    (P �``��       (8Pp��`���         �@�@X '   @���Xx'?                                         p               ��   ?k?ag44  ??__,?,?      � ��� �  �      �������� �                0�(�l�D����<<   p�8���������<<                            � �             � �              ~      ~      ~      ~      <   <          <   <                                   	 : x 0   		::xx00     
 
 8 8       



8888                             @              @         @@��ND         @@� N (8 .; ??;;� � `����0�\�� ��@�������|��܈�    ` �`h04~�L    ``��xx<<z~���nz4h0�``     ��~~<<xx��``     (>}�x| 88>>��|| $ 44444 <<,<,<,<,<,< (>}�x| 88>>��||    ~ � �|~         ~~����~~      ww�o�Q�a�x�  w����������      ����������      ����������            �� �P�(�t��    ������������        !?Ro        ??o (P �@@�����(8Pp��@�����  :=1>2=5:  =?>?=?:?������ ��p|�� � ��������p��� � �5:s|uzr}9>:?|z}>?   �@����D���  ������D�����    @ �@Q!)    @@��Qq)9  88||�������\�  88||����������    !;E4K   ?!?EK  ��@��` �0��p�  ����`���������4K:E4K%    KEK%?    p�p�p�`�����    ������������    � ��      �����      �������!�sz�xx  ������������xx  :G>A"!   GA"?!?  8��|^��^�>�\�`���|���^�>�\�����2=        =?        �0�P(�((((( �h���(8(8(8(8(8
( 
(8<���`� `        ������``        	
        ��<�8ĸD��0��  ��������������  :Ŕ��G>>  ������>>  ���Д�
     ������
                          x � rp���|x��  xx����:�����8�< N�>�.�Fn,,<<r~������r~4<4<                                     ,,,,,    4<4<4<4<4< 2����>> .>�������">        < N��&        <<r~����             ���             @���            ,,,,,     4<4<4<4<4<                                    n���N~<<     r~������B~<<           ?         ?? ?    w.,,,,   y2>4<4<4<4<    �  � x�8��@� � �����������H�H�  � � � � � � �   H�H�H�x�@�@���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  � � � � � � � �  ���������  ����� ���������������    /         ??????    ������    �����������                   ���0�0�0      ���������                                @�@�@          ������� � � ����� ���x�p�`� � ������������ ��������� � � ''/ ??     ???? ? ?    ���������     ����� � �                   �0�������       �� � � � �                            �����            � � �          ��<�x�x�x�<��             �<�x�x�x�<���            ��~�$~���:��t�N� � � � � � � ~ � <��� � � � � � �  �    �   � �f~�� � �� �   g �   � < � 8 �"��4��}'��c�<~�3 � � � � � � � 8�8��?�x�������           � �8�x���8����     0       ��p�����<�0�              ��������p�0�            �����{�|����� � � � � � � � ���~������� � � � � � � � ?�a�� ������� � � � � � � � ��{^���~����� � � � � � � � � �$$�Z�~�<g�>� � � � � � � � �3�9�\�.�.�\�8�1 ?  � �  ?  ����������?        ��@�?��O�9���  ?       @   ��@��?�?�?�?�?  ?       �?�� �@���~�   ?       � � ����0��� � � � | ~ ~ ~ �
��X�0�� � � ~ ~ ~ ~ �    � � ��(8������ �D�    � 8 | | � � �_�_�~�p�~�_�_�_# / ? ? ? / #   ���a�a�a�a�a�~ ~        � >?>?AA���  � � � � � �   � �`�`�`��|�~�~~           � |w|w�����   � � � � � �   � � ��J��_���       @ @     � ��/�Z�\�W�S�Q� � ` A A @ D F �P�X�\�_�O� �� A @ @ @ ` p � � � �O��9�s�g�N�}         8�x�����������x�   @ � � � @   `�������������x�          � @   ��~�>����w��� � � � � � � ~ � � � ��� � �  � ? � � 8  � � � �f~�� � v�� �   w �   � �   �J��U����;o���~k � � � � � � � ��x�?�<�8�0�0��             ����x�0��8�x�              ������������       @ �   ����������P             ������7��8���� � � � � � � � ���~������� � � � � � � � ?�a�� �����z�|� � � � � � � � ��{^�?�a������� � � � � � � � � �$f�>�\�~�>c� f � � � � � � �9��n�7�7�g��8?   � �   ? ����������?        ��@�?��O�9���  ?       @   ��@��?�?�?�?�>  ?       �>�� �@���~�   ?       � � ��$�F�H��� � � � ~ ~ ~ ~ ���T�j��� � ~ ~ ~ ~ �    � ���D|������ �D� 8 � | | � � � �_��|���|��_�_' ?  �  ? '   ��������~ ~ ~ ~ ~ ~ ~   �  AAAA���  � � � � � �   � � � �@�>�`�p�|~ ~ ~ >      � ����	�	��   � � � � � �   �� � �
�N�_���       @     � �� �G�O�Z�\�W� � x ` @ A A @ �S�Q�P�X�L� �� D F A @ ` p � � � �?�s�g�F�^�}�s         ����������������            ����������������      � @ ��|�<�)}����V�,� � � � � � � � � � � � � � <��� �  �   � �  � � � �f~�� � f�� �   � �   � � �R�������b�>~��f� � � � � � � � p�������`�0�<��  @ �         ���������              8�0�0�8��?�s���            ���������0�         `   ����7��8���� � � � � � � � ���������� � � � � � � � �0�p�������z��� � � � � � � � �}���p������� � � � � � � � � �B�f�<~�<Á~C� f � � � � � � ��f�3���3�f�?   � �   ? ����������?        ��@�?��O�9���  ?       @   ��@������  ?       ��� �@����   ?       � � ��0�`�@�b�b� � � � ~ ~ ~ ~ �B�@�d��� � � ~ ~ ~ ~ �    � � ��  ������ �D�    � 8 | | � � �_�_�^�^�^�_�_�_# / ? ? ? / #   ���y�q�q�q�q�~ ~        � >?>?>?!!���  � � � � � �   � �p�x�|��~�~�~~            � |w|w|w�7���   � � � � � �   � ��@�
��_���     D @ @     � �� �@�@�G�O�Z� �  p ` @ @ A �\�W�S�Q�@� �� A @ D F a p � � � ��g�N�]�{�w�n            $ N��>��  <<r~��������   <~ ���$�$  $<B~��������   ,Z�8�4�d�l  4<f~���������,�>��vn,<   ��������R~$<  �$���N<   ��������r~$<  �t�d�h�X~ <    ��������B~$<  � �g�g�g�g�g�g�g� � � � � � � � � �������������� � � � � � � � �`�`�`�`�`�p�� � � � � � � � � �������� � � � �  � � � � �`�g�g�g�g�g�g� � � � � � � � � ��������������  � � � � � � �g�`�`�`�`��� � � � � � � � � ���������� � � � �  � � � � ��`�g�g�g�g�g� � � � � � � � � �������������� �  � � � � � �g�g�`�`�`��� � � � � � � � � ����������� � � � �  � � � � ���`�o�o�o�o� � � � � � � � � �������������� � � � � � � � �o�o�o�o�`��� � � � � � � � � �������������� � � � � � � � �   < F8/   ; )   < z 1   , >  2l � � � � �  . T � � � � ^       @ �@�@_ ;       @ � � a $       � � � �      y � � � ^             ?             (         8 � � �         8 � � �    w+T+T+ \#U+   w w w T w w   � ��*�*�� :�j�  � � � � * � �    w+T+T+ \#U+   w w w T w w   � ��*�*�� :�j�  � � � � * � �  =3=13   > ? > > ? � �@�0�H�0�H�p�8� p � | � | | �  =3=13   > ? > > ? � �@�0�H�0�H�p�8� p � | � | | � D " 1 Y o � o       q Z F b 2    ��� �<�>�   �  � �  ?   	             ���=�&n     ~ >  � � n       	             ���=�&n     ~ >  � � n     / ~ �@�@\ 3 < q � � o 3   � ���=�&~   _ ~ >  � � ~   w+w*A> w*w+@? w w @ ~ w w @  ���T�|� �T���� � �  ~ � �  � w+w*A> w*w+@? w w @ ~ w w @  ���T�|� �T���� � �  ~ � �  � ?<8 ? ? ? ? ? ?   ? ?   ? ��<���� ���� � � �  � �  � ?<8 ? ? ? ? ? ?   ? ?   ? ��<���� ���� � � �  � �  � '  < i * 8  / _ >    �n  �n�� � �  � � � � � � �         ?	       
   5       ` � �@� ��      ` � �  �        	       	          � ����80      �   H �        ??       	  ( 2       � ��������      �   P P                        	          � �@�@ܠ        0 h � d                      
         p �@�@�         p h h �     ` � �}"ZY    ` � � W m j      ? O0�@]��f     9 u � � Y       < zU*$%      < F { ; :       < Z$�hj��T      < f � � Z                                                                 __o!~z |47 r w X k _ K 6  �0���~^>,쀀 N �  � � � l � >?/o/k+; !   0 P T $   |x��������\Hx`� �   & " � � � ?/ * 0 $   ; ? /   ���@h h ��8��� ( � � � T � h � /.37   9 7 < 8    � O��Z�l�p8�� � � u � ~ | � � � ".5
&>   ; ? ; 9 9   ��쐖hV��44�� � d t � � > � � � ��C<;<   | s } < ?    7�{���p<�� � � . � � | � � � � M2�f�fa8   r � � ~ ?    �H�$�,�$<�� � � L & . > � � � �                                                                   f �f�~�f�f�~r<  ff����������~~      ` �@�`�pz8      ``�����F~44<2<2< <<<<<<>><<>><<99z8�p�`�@`   '?'?F~������``  � �������                � �~�}�{��?�\�l       ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���� 0 	  	  
  
  $   ����                �x        �          �                                                                                            D J                �       !'-39<BHLRX]ciouy����������                               $(,39=DGJMQW]ahnsz~��������                                 &,06<AGMSVY^dkou{��������                                        !GIR  ��V     �    ��    �i�    ��9    � =C     8�   �    c��!s>9WN��c��!s>9WN�  �k-�R�w2%��%�c�-�+�  c����M}{�c��	�+�  c�0*���$�c�S)Bc+�  ���5�s)5��Y�c��	�R�s  c��&)}���c�  ��  �=;�fR�B)&�Yc��!s>9WN�  ���J�?�  �y��9��f�E  �Ii�b�o�QO~  �Z�U�v��*�  ����6��A%  �������  ��1��6�V~�e  ��IS;�_7  �~#u�6�q`  ��'-^��z�d  ��2� >&��V�9  �k-�)�/%�w�R  �~#��6��x�YG6h;J
�\*qz  ��V     �    ��    �i�    ��9    � =C     8�   �    c��!s>9WN��c��!s>9WN�  �k-�R�w2%��%�c�-�+�  c����M}{�c��	�+�  c�0*���$�c�S)Bc+�  ���5�s)5��Y�c��	�R�s  c��&)}���c�  ��  �=;�fR�B)&�Yc��!s>9WN�  ���J�?�  �y��9��f�E  �Ii�b�o�QO~  �Z�U�v��*�  ����6��A%  �������  ��1��6�V~�e  ��IS;�_7  �~#u�6�q`  ��'-^��z�d  ��2� >&��V�9  �k-�)�/%�w�R  �~#��6��x�YG6h;J
�\*qz  P(V�R([([(\( �<  �,�, � �  q(   �(�(�$�$�h�h      T(�<X(�,�,](�$�$�$ �$�$ �$�$ �$ �$�$�$           T(�<X(�,�,](                          T(N<Y([�[�\�                 %%       T(^<Th                    %%       P�V(P�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����������������� � � � � � � � ����������������� � � � � � � � ����������������� � � � � � � �                                                                                                                                                                                                       � � � ��              �                                                                                                                                                               ???�?����   ? ?   � ����������������� � � � � � � � ����������������� � � � � � � � ����������������� � � � � � � �       � � � ����            � �                                                                                                                                           ����������������� � � � � � � �                                                                                                                                                        ������� �       � � �           ������� �       � � �           ������� �       � � �           ������� �       � � �           ������� �       � � �                                                                                                                                         ???�?����   ? ?   � ����������������� � � � � � � �       � � � ����            � �                                                                                                                                                                                                                                                                                                                                                                                                ��                              �                                                                                                                    ��                          <                                                                                                                                                                                                                                                                        � �                                                                                                                                                                                                                                                                                                                                            A A    @ @  @          �                                                                                            � � � � � �U                              ��                                                                                                                                                                                                                                                       �l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         :>� �6c *� � �V� �V4 "W4 *W4 &X4 &YT *HT JHT *Tf <8 ^F, (* (B R[ G$GII$IJ J ^X� �� X� �� �� T� $T� J� $J� K� $K� L� $L&hX RZ� �J ^Z `WK `I� "E� �D� K� "K� �J� �K� �K� �LF $� � } 8	� ^� `Z� dW� `� �
� Wk � I� T� �
�  W� $X� Y�  Y: `N<X@X4Z8Z<ZDZHZ@[D[� U� $U� V� $V&`T&hT&\U&`X&lU&`V&hV&pV&\WM �[M �[M �\C ���	�	��� ������ �����  ʌ���t ����� prpL��! ������" ����S �hd��s ���� (Td��2 ��C ���	�	��� ������ �����  ʌ���t ����� prpL��! ������" ����S �hd��s ���� (Td��2 �����B ����� (��j ����� ��$��� 
$��U P��A >p���I \��p��� PlPl��� 2	J	�����  2 ������� 00��� 00��� P��� h��= LpPl��2  � �    �    xx�      2 �                                                                                                &&&&
  
                                                                                  * ((**   (
 (*                              bb  $$          bb'''    $    '''''   $    '''''$    ''''' #   ''''' 'T  ''''''''T  '  "        						'' '``  Kggggffff        'c'UUD  :; 'c'SSD   				��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �                                     � �             �            P l{4          p | w          
6�,          > �      337       ? ? ?     � ��~D;����    � 4 � � g     
              � �`��,�p_��  � � v r � � �    >     ? O K X   � ��0�<���� ��  � � � � � � : ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �                  � ����x|8|8|   � � � � | | |   �c�h�	��n} � � � � �    =���� �l�r�|| � ? ?  � � � | 7?   ? ?        � ����0p�� 0 � m " b � � � 0 3?/&    ? ? 3 :  ���l���`� �     � � � � � �     ��A�dw	> � � � z /    ���^ |0 � � } � � � � � �    /7s      ; , O   � ��0�8�����0  � � � � � 4 �    ?7       # *   � `�x������8�p  � � � � � � r           P l�t          p | �          
6�.          > �           0 H0w          0 x           
�           �             8 '            8 ?            4�0           < �             8 '            8 ?            4�0           < �  0g8�p�`� �                � ��������             �8�?�8�;�;�;��            �4�����������       � � � �   ���`0? � � � H 6    �y�����p��� � � 	  l � 0 � 3?77]8 - 8 / , z '   � � � | ���p��� � � � � d � 0 � �c�(�I�L}- � � � �  ?   =��m��4�x�x�pp � ? ? { � � � p �s�@�{7< � � � O ?    <���<
�4����� � > � � � � � � K5V)v	[$j4; G O o   ?   ��x�x��z\�0�� � � � � � � � � M3Y'w7/	 G O  ; 9    � ���t��ĸ�0�� � � � � � � � � �9�
�e�b�a�p�8�8              ��y��C�`^�*ՙf�7               W/X'_ [$K4c0                 ���������                <6>}"    ? ? ? ~ � ��� �0��(�8�� � � x < l | >  8 ; lE:L7, ( + _ _ ~  ?     � r̹n�.�v�    � �  ?  �  :~      ?  � @��@� ��(�|�.؀ � � � � � � �    /s,]n)     1 ]  W ~ �B�������~��~�~ � � � � � � �      /3}"       1 = _   ~ �B�������~��  ~ � � � � � �     � ������0�D    � � � � � �       /3        1 =   ~ �B�������~��  ~ � � � � � �        , < $ 4        4 < < ,         ` � ��        ` � � �            ��(           � < ^#! 7   { y >    z������X0�� � � � � | � p � ??_ 0w(: ? ? s O _ ?   .�����,�p|���� � � � � | � � � _/.~=<    ?     ���t~�<����0�@� � � � � � � � � 17    K ;        $����ý�<~�<�� � � � � � ~ < � ^o)?  g W +      ~�$�����=g��X� � � � � �  � � z�����@Ȱ� �   � � � � � � �   =o-/';: / S 3 ;  ' &  ~�$����ý�<�� � � � � � �  � 444 $        , , , <        ?_%L0~ ?  ? ~  s 2    <�������@� 0�� � � > ~ � � 0 �         ` � ��        ` � � �            ��(           � <         @ � ��         @ � � �           p �0�P          p � x      ={$_O	      # ] g w         ~ �~��<�        ~ � � �        ={$_        # ] g           ~ �~��          ~ � �       0 X �@�$�      0 h � � � 8 < z4][O /	  < N k m  7        p �p�~?���      p � � � �  8  T T |                        D � D                          < f$�B� �       < Z � � �  8 llllll ( T T T T T T     ?  �? ?       ? @ � @ ?   ?_%L0~ ?    ? ~  s 2     <�������@��p� � � > ~ � � � � ���~}3{A>> � � �   { A > x��h�X~������   � � � � � � �   /	    7         �����<~��~�<<�� � � � � � � < � O	/	    w 7        <������;{�ƽ�? � � � � � � � ? ����@P��  �� � � � � � �   � �                    ���?�α�= � � � � �    8 (((((((8 ( ( ( ( ( ( (       � ��           � � �     �$��Z $      � � � f <      | T(D8(| D8( D l | 8 | D (      � �d�6�d�       � z 9 z �        /?^#_1      7 7  {      (�0��z���     8 � � � �        /        7          (�0��x�       8 � � �    /    7        (�0��p�����   8 � � � � �  / 7 ?      ?     � ���������    � � � � � �      =6        ?      � � � ����m8    � � � �  �      =6        ?      � �`�0����}8    � � � �  �    //7    >   ? /       � p�8��(��      � � � � �   ??~7     ? ; w � ��� `���� ���� � � � � � � � �m�C��K     � � � � O 
    ������u@� p     � � � � � P     ?''36 ; = ? ? ?    �����̸l8�0x0 � � � � � � x 0 73   ? ?        ��̸�p�p�0p     � � � � � p     ;7	 7 ?       �0��x��������� � � � � � � � � '�o�~     w � �        �<�|�������     � � � � � �     '�o�~       w � �         �<�~���88       � � � � 8       .?	?	?   ? ; 9 -      t������������   � � � � � � �   |??      ?        �x������ݸ�t`� � � � � � � � �                                                                   ??~7     ? ; w � ��� `���� ���� � � � � � � �   7'      ; 9   � � ��:�~���  � � � � � � �  .'/    ? ? ?  � ��p�8�t����xx�� � � � � � � �  ?2�c�g|?~  ?  � �       � � @�@�@��     � � � � � �  ?13>?   ? y s ? ?   � ���  � � �@�  � � � � � � �    <x���    3 W � � �   � ��|0�O    � 0 � 
 � � �       ` �`�`�@      ` � � �         ���         � �                                                                 |??      ?        �x�|�����8�t`� � � � � � � � � /.   = ?       ��t���� p@� � � � � � � � � ` � 7      ?   x�p���8�p�� ��� � � � � � � � � O~? _  O  w '   � ����m����   � � � � � �    ??'> /  ' ? ;    � |8n<�t��5���� � | ~ � � � � � �w5:;  � J / $     �T �����  � Z � d   �  n=n;>8       ? 8       v�v�<����       � � < � �       �m�a�]�>����]e�A��>����]����k��x�i��6�V������r�`��T��`�s�_�o�?e>	w,`�3�W�O�'�	?$    ? ??=;?     ??????@ � x > =   	 @@��Xx&>#?    � �0�:�y��  ����������  c �  ?    �?? � �f�B�f�<� � �  �f�J�f������� �  ( ( h h h �   880x0x0xp�  4 : z z } �  <><~<~>~�  8??????  88????????????      ����������      ����������                                ����            ����1111! !//????? ? ? ?L L L L � ���xt8���������� � ����I�I�+�^�c��� I�I�*�\�@��� ��X_���?����� P�B�
������� �    ���  ���        �� �����     ??� ??�? {???G??����?�����o��y�����������������      ? � >          ??�?       � ~<= � �        ������� �� � ����� � p�`�P�P�P�P�`�p�� ������� p�n�Z�P�T�Z�n�p�????1     ????????1?     �����������<� ����������<��               �����������     ���������� �    /�_� �@  ?    ��?� �8� � ~ ��� �� ������������� ������������������������������<<B~�ý��[g~Z$$<<~~������gZ~$$�$�$�$�$�$�$�$�$Z�Z�Z�Z�Z�Z�Z�Z�,,vF����nn<< <~\�8�~ <  204z   ???E� ��8 <0< �� � �����������B�ǂ�B@?@?�?����?��B�" ������A�B��������A�B�D�H� ������� 8?8???????????????� �����<����x�8����������������                       ������          ������               ? �;����������  ??������� �?�?�?�?��!^�� ���@�H�^�!� � �� � ���䅄{�  �������z��� �������������������������������$�$�$�$�<�~ < Z�Z�Z�Z�B�f�<~ <8 D8�|��f~,<  88||��f�,~< 4,4,4,4,4,4,4,4,,<,<,<,<,<,<,<,<��Lo0 ~?  ����{~S/?����� ~�� x�� �����~������������@?@?@?�_������ "B������������A�@���� ��D�B�A�@�?=???> ????????????�8�x�x�x�xl���� ����������������              �����������00   ����������0� 0  ???x8`  k6k6 ? ?@G_ww������
����������@ @ @            @ @ @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (((((((((((((((((((((((((((((((((          ���������� ��U� � � � �0� � � �� � � �� �0������'?���;�}��������������?��~w�n������ � �`����������������������f���� ���?�^������ ����_��)�;��s� � � � �@������� � � � ��o���x� ��
�
�
��{�[�0�/�_�_�w��(_��y9�� �w����;���3������u���� � � � � � � � ������������������������������>�������������������MZ��_Y�~��������������������������������5�m��~���V�g���������y��|~� ��3_�����?N����w����د�c��������������G���[�S�Q�Y�$��c��7�/�_��������t��������F������7���������{}�����W���E� ��UU�����U���T� ��UU�� � � ������ �`W��x؏�������]���������}��n���������������������������+���������������������	������m�g�������(�S��?�����������g�� ����A��������7���w�����;��8�<_������|�8����{�������O�7�}��{��������0�������������������e�������������������g�c���{��������^���W�� � � � ���?�~��?�?�?�?���������������+�����������������8�������y��������<�x���c���������9������>��<�<���?���o�O��N&��L����ȿ�������� ���g=�<���	� � �o��z������ <� �������?��������ܿľǇ������s:���v�=�s���� �������{���������o������}:�������������+��?��'�_���������������������ӯ�ϳ7�G�V������ � � � � � � � ������� � � � � � � � ��� � � � � � � � ����� � �@�@� � � � � ���� � � � � � � �  ��?������������s�o�~�p����������� � � ����?h� � ������>�c��<�x�xw�w�y���r���������\�����������������n������ � �����p�0�;�� � � � ���@���?����� � � ������ � � �� � �@������ � �����+���� � � � �8�� � o��`��p�>�ͳ��2�������������������b������������?���O�F����g�;��~�g4�d����������������X���������������������l�(������������5��?N�!�?�<���x���?��?�� � � � � ����� � � � � �>���|� ��������G�z��>����{���'�'��_�����߿�� � � � �`�0���`?��� ��� � ������������������������������`�p�?���?g�3�t�i�����������~�������������B�F������o�O�l�*߷K�����ü����g�X��^��>�~m�����o� ��h�H�M�G�a�1c�8�~����]�]�����~�����������W�_�_�_�\�Y�Y�;��g����������}�=���������2������`��� � �?���p�8�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��	�������	����																																																	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
					
	           
                  	                                   
        
											 		   	� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � X�N�F�@�:�4�.�*�$�"�����
���� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����K�g�������������������ہ�S������]������������������j���:�������_���،������:�k�ڏ����������ݔ����ș	�6�L�j���Ț���D�k�y������A�~�Ȝ�q���ڝ�P�|����&�a����1����)�j����*�f����_����7�������?������(�q����,�a�����K����'���'�����$����������-���ޮ�9�u���ݯ�4������O����������o�����^��X��q��<�v�w���ߺ�=�K�f�y���Ի���i����ν��e�ؾd�����D�����7����O�����M������@�h������,�]�%�~�����*�o�����!�N�v������F���v������������>��D�~�����(�k�����)������K������L�����
�i���)�����X��?�Q���-�b��������@���_���R������[������������`����� �8�L�o����[������?�z�����+�c���v���Q���g���x���������=��P���;��� �����@����������	�/�c���+�:�G�b�~��������J�3�^�T������Y�{������@�p�����"�Y�w���������p���O�g���'�c������1�[�#�������.�����W�r��m�������!�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��V     �    ��    �i�    ��9    � =C     8�   �    c�,*=�Itb���c�,*=�Itb-�  �k-�R�w/%��)�c&-�9�=&-*=-  c�,*=�Itb���c�$)G1�$�,�  ��%�!������
L!56K�o  �!�5�sA��a�c�$&-�9�9sN�^  ceIiQ�Di]O~�c�(�$���I*=  �=;�fR�B)&�Yc�,*=�Itb��  ���J�?�  �y��9��f�E  �Ii�b�o�QO~  �Z�U�v��*�  ����6��A%  �������  ��1��6�V~�e  ��IS;�_7  �~#u�6�q`  ��'-^��z�d  ��2� >&��V�9  �k-�)�/%�w�R  �~#��6��x�YG6h;J
�\*qz                                  �                               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           l                               	                                  @A                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       |Y0�                P                 `          � 3 w �  3                    3         ��~  �����        ��~  �����        ��~  �����        @�~  �����        ��~  �����   �����������       &�� �� �� �       &�� � ��  
�          J  X}76                    3    ll            �   ��G(          T  �         T       8��      d          =  � %           ���             �             �                    �                      �  p `      
              �                          @   	                           <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<������������������,�-�<<<<<<<<<<<<��������������������������������������<<<<<<<<<<<<���������������������������������������<<<<<<<<<<<<����������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�������������������������H<<<<<<<������������������������H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<�����������������������H�H�H<<<<<<<-�,����������������������H�H�H<<<<<<<���������������������������������������������șH�H<<<<<<<�����������������������������������������������ȒH<<<<<<<��������������������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<����������(�(<<<<<<<<<<<<<<<<<<<<<����������(�(<<<<<<<<<<<<<<<<<<<<<����������(�(<<<<<<<<<<<<<<<<<<<<<���������,(-(<<<<<<<<<<<<<<<<<<<<<�����������<<<<<<<<<<<<<<<<<<<<<�����������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<��������������������<<<<<<<<<<<<����������������������<<<<<<<<<<<<��������������������������������������<<<<<<<<<<<<���������������������������������������<<<<<<<<<<<<����������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�(�(���������H<<<<<<<<<<<<<<<<<<<<<�(�(��������H�H<<<<<<<<<<<<<<<<<<<<<�(�(�������H�H�H<<<<<<<<<<<<<<<<<<<<<-h,h�������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H<<<<<<<<<<<<<<<<<<<<<���������H�H�H���������H<<<<<<<<<<<<���������H�H���������H�H<<<<<<<<<<<<���������H���������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<������������������H�H�H<<<<<<<<<<<<�Ȱ�����������������H�H�H<<<<<<<<<<<<�����������������������������������șH�H<<<<<<<<<<<<�������������������������������������ȒH<<<<<<<<<<<<����������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FPQPPQPQPQPQPQPQP���������������CGa``a`a`a`a`a`a`���������������STHpppppppppppppp���������������CDq��P��P��P��P��P��P��P���������������CDq������������������������������STq�����������������������������CDq������������������������������STq�����������������������������CDq������������������������������STq����((M�����������������������CDq�����88M�����������������������STq�����������������������������CDq������������������������������STq����((M�����������������������CDq�����88M�����������������������STq�����������������������������STq���Ь��Ь��Ь��Ь��Ь��Ь������������������CDH�p�p�p�p�p�p�p�p�p�p�p�p��x����������������SG�a�`�`�a�`�a�`�a�`�a�`�a�`���	���������������F�P�Q�P�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������8�8�8�8�8�����������������QPQPQPQPQPQ(P(Q(P(�(�(�h�hQ(PQFH����������a`a`a`a`a`a(`(a(`((�	�	ha`GHCH����������ppppppppppp(p(p(p((HpHHTHSH������������P��P��P��P��P��P��P��P��P�PqHDHCH������������������������������qHDHCH������������������((M���������PqHTHSH������������������88M����������qHDHCH�����������������������������PqHTHSH������������������������������qHDHCH������������������((M���������PqHTHSH������������������88M����������qHDHCH�����������������������������PqHTHSH������������������������������qHDHCH�����������������������������PqHTHSH������������������������������qHDHCH�����������������������������PqHTHSH�������������Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ь��Ю�qHTHSH����������x��p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�H�DHCH�����������	�a�`�a�`�a�`�a�`�a�`�a�`�a�`�a�`�a�`�G�SH����������Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�F������������L�H�H�H�����������������������������̥H�H�H�����������������������������L�H�H�H�����������������������������̥H�H�H�����������������������������L�H�H�H����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FPQPPQPQ������������������������CGa``a�	������������������������STHpppx������������������������CDq��P��P�������������������������CDq������������������������������STq��������������������FPQPPQPQPVTq��������������������CGa``a`a`aWq���������������������STHppppppppX��������������������CDq��P��P��P��P���������������������CDq������������������������������STq�����������������������������CDq������������������������������STq�����������������������������CDq������������������������������STq�����������������������������STq���Ь��Ь��Ь��Ь��Ь��Ь������������������CDH�p�p�p�p�p�p�p�p�p�p�p�p��5����������������SG�a�`�`�a�`�a�`�a�`�a�`�a�`�$�%����������������F�P�Q�P�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P��������������������������������������������������������������������������������������������������������������������������������������������������������������������̥H�H�H�����������������������������L�H�H�H�����������������������������̥H�H�H�����������������������������L�H�H�H�����������������������������̥H�H�H�����������������������������L�H�H�H�����������������������������̥H�H�H����������������������������PQPQQPQFH�������������������������	H`aa`GHCH������������������������xHHpppHHTHSH�������������������������P��P��PqHDHCH������������������������������qHDHCH�����������������������������PqHTHSH�����������������������������PqHTHVHPQPQPQPQFH���������������������qHWH``a`a`a`GHCH��������������������PXHppppppppHHTHSH��������������������P�P��P�P��P��P�PqHDHCH������������������������������qHDHCH�����������������������������PqHTHSH������������������������������qHDHCH�����������������������������PqHTHSH������������������������������qHDHCH�����������������������������PqHTHSH������������������Ь��Ь��Ь��Ь��Ь��Ь���qHTHSH���������������5��p�p�p�p�p�p�p�p�p�p�p�p�H�DHCH���������������%�$�a�`�a�`�a�`�a�`�a�`�a�a�`�G�SH���������������Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�Q�P�Q�F�����������������L�H�H�H�����������������������������̥H�H�H�����������������������������L�H�H�H�����������������������������̥H�H�H������������������������������������������������������������� �`�o�o_�m�}��7`�� �	��7����  ���}G<<YB�� ��� ���������X��  ����#�#�$�)� ��� �������������p�{��0�?�?�? ������P�O�O�_���7�������O��� � � � �"��������?�?�?�?�>�<� �<_�_�_�_�^�]�B��O�G���G��B�
���������,���p��� � �  ���  ��  � � � � ��� � ���x�x�xC�c�s��<`� � � � �0� � ���p�{�{��� �  ������ � � � ���7����� �� �  � � � �"� � � �}��$��>������� ���
� �}��&��>���� � �� � ��� �s��#��;���� � �� � � �� �~��'��?����������
� �s��#��;���� � �� � � �� �}�o�$�<��������� ���
� ��P�3I��� �Z� (�����6�b�B�� �+��� �������� ����������� � �    ??11##''..<<  @@q@c@g@n@| � ���?�?�?�� ��a�`�@�@�@�`� � �� � �@�� �������������������� ���   �� � � � � � ��� ���� �?� �?�?�  � �� � � � �?�s�c�#�;������ � �� � � �� ��1�;�w�n3�l��C�? � � � � ��� �?��u��>?������ � ��0��� � � �U��*�������O��� � � � �"�������U��*�������y��� � � � �"� � ��U��*����� �� �  � � � �"� � � �U��*���������}~ � � � �"�������U��*����� �� �  � � � �"� � � �� �o�o�oZ�j�z��7`�����7���� ������������_` �����������������p�{��p��� ������ ������7���������}~ � � � �"�������� �o�o�oU�m�}��7`� � � � �0� � ��  ����?���� � � � � � ���`���p�{��x��� ������ � � � ���7�������y��� � � � �"� � ��� �o�o�o\�i���4`� � � ��2� � ��  �~�<~���Z�$� � � ���B�$�� ���p�{��p��z�t ������ � �����7����� �� �  � � � �"� � � ��  � �� ��=�}�  � � � �y�@� � ��  � �� ����  � � � ��� � � �� �������> � � � � � � � ��4������a�� � � � � � � � �~�m�'�?������������
� �����Z�P��@���@������� � � � ��~�}�� � � � � �~� � � � � � ��������_�?�_�?p��� � � � � � �}�j�&�>������ � �� � ��� ��������I]��� � � �A����� ��a�`�p�x�|�~����� � � � � �������szy|sz���������������{�k�#�;������ � �� � � �� �� U��U � � ����� � � � � � � � ��h�t�z�}�}�z�t�h���������_�?�_�?�_�?�_�? � � � � � � � ��h�f�f�f�f�f�h�f ������ ���f�f�f�f�h�f�f�f���� ������p��� ������ �p�� � � � � �f������� ���� � � ���� � � �    ���̄�  �����8800  !!##??    @x@p@`@a@c@  $$DD����    &F����  �m�m�m�m�l�m�m� � � � � � � � �U�U�U�]��*U�U�U� � � � � � � � �f � �     � �    f � �     � �  � �?�_�`�g�k�l�l � � � � � � � ���`�_�X�W�V�U� � � � � � � � ���d�_�Z�w�^�U� � � � � � � � ����nr�d��v��,�I� � � � � � � � ��l&�M��6�m�� �I � � � � � � � ���$�I}��$�Im��% � � � � � � � ��?�~� �B�~�~�~�~ � �~�<� � � � �� � � � � �B�~�~ �~�~�~�~�<� � �� F�B�)�`���� ��=�V��y�m��� �?� )�`���� � � �V��y�m���  � �� ���  � � � � � � � � �� ���  � �� � � � � � � � � �        �m�m�m�l�m�m�m�a � � � � � � � �W�U�U��"U�U�U�w� � � � � � � � �" 
 �  b   �    " 
 �  b   �  m������ ���@� � ��� ��W(�jU�����|��� � � �� �� �]"�h���R�U�� �� � � �� � � �� � ��H��K�5�{ � � � � � � � �����+��	��- � � � � � � � ��������g��n� � � � � � � � �            �                ����~�~�~�~�~�>�>�> � � � � � � � �?� �� J��a��� � � �5�w��� ��  ���~���{�  � � � � � � ��� � �� �� �� ��  � � � � � � � ���  �� �� ��  � � � � � � � �<�~����������|� ���B�$�����|�����������<������ ��$�B�� ������� � � � � �!�!� �ww����-��>������@��� � � �����<���� � � � � � � � �>?:;tw���\��� ������� � � � �� ��� ��� �  � � � � � � � ��l�l�l�`�l�l�l� � � � � � � � ��� �< �   �   � � � < �   �  0��@�H��"@� �� � � � � � � � �  (���  (���    � � � " � � ��>�>�>�>�>�>�� � � � � � � � �� 7�m� � �� �� � � �� � � � ��� ���� ��  � � � � �� � � �� �� �� ��  � � � � � � � �W�U�U��"U�U�U�w� � � � � � � � �Y�,s<3^9^9�s�wX� ������������� �C���z�:ǋ����Ӡ� � � � �@� � �ms|st{���؍���������P� �@� � �78���������� � � � ��� ���������g�c��� �@� � � ��(�5>�����د�������� �� �@� � �� U��U � � ����� � � � � � � � ��_�?�_�?�_�?�_�? � � � � � � � ��B  �   �       �   �   �     @?� � �� � �(�  � � � � � � � �@*�(�
$�  � j � : �  � ��������  � � � � � � � �� �� ���@�� � � � � �?� � ��=�7� �?� ���  � �?� � � � � �    5k������������������]<�ys����ϟ�??�������0�`���� �   � s�� �B������� ���0�c�� �   � v����m�������� � � � �m��������� ����������������������������������������� �   �  ������������� � � � � �� �   �  ������c������ � � � � �� �   � �}��� ������ � �}�}� �� �   � � � ������ � ����� �� �����������������������������������������������  A~�~�~����������� � � ���@��߿߿߿o���?� � � � � � ������0���� �� � �� � ���|s���� ��0�0�G��� � � ��� �� �   �  ������������� � � � � �� �   �  ������������� � � � � �������������������������������������������������� � � � ������������������������������������ ���� �  @ ?�?�?�?�� �����@�@�@�@� � �    ���������� ����� � � � � � �>?>?>?>?>?>?>?>?����������������>?>?>?>?>?>?B ?����������������~��~���������� ���B�$��� �@���ls�g��s��?�w� � � � ��� ���@��(�A�#�C�	� � � � ��� ���� �����  � �������������    //+75;:=<?����������������>?>?��������������� ����� �������������������������������������������������   � � �� ����� � � � � � � ��� ��?�� �� � ��@�@� � � � � �wwwwww����������������� �wwwwww
st����������������  @? _opwuv�����������������wL�,��������� � � � �� � ����������������������������������� � � � � � � �wwwL�����`������ � � � ����>�|v������o��>�|����������� �� � ���������  � ����������� ��>�>�>�>� �>�>�>>�>�>�>� �>�>�>�� � �?�?�?�?�?�> � �?�?�?�?�?�>��>�>��������� >�>����������� �� ���	3�g��B� ������0�c�� �   � v����m�� ����� � � � �m��l�j�d�h�Q�!�B� ������1�a���������`�a�a�`�a�a�`�a�� �   �  ������������ � � � � ��  �O���'� � � ��0�c�G�@�� ��  � �����  � ��������������� �����  � ��������������� �ȟ�/� � � ����0�g�O�@�� ��  � �����  � �������������  ������������������� � �>?>?>?>?/0 2���������������0� ?~?>?>?>?>?>?GF������������������_`#<=>>?>?>?>? ���������������wsqpc0���W����������� � ���Lw���s�5x<Gw@��� � �������� � � � � � � � � � � � � � � � �                                 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ������������ ����������� � � � � � � ����� � � � � � � � �� � � � � � � � ����������������� � � �  7 M � ������������������6�{rͺ�K�������{�����������
�)� ���� � ���������������� �<�<� �=������<�B�B�=���$��!�>�� � ��������A�b��������                                                                                                                                �������������� ��������������� � � � � � � � � � � � � � � � � �                                                                                                                                                                                                �<�v�2�2�^�X�p�P��v�2�2�^�Y�s�W�� �B��0���� ������;��������� !�?�?�?�� � ���!�@�@�@�!�>� �`d � sm^��ޛ�p�������!�!�!�                                                                                                                                                                �&� � �<� �~�~� X�Z�B�B�~� � � �� �`��?�?���  ���@�@� � � ��B�$�f�f�f�f�f�~������� �� 	w��ϼۼ[�[� ��������������[�I�d�0ϼ����������������������@������V�V�F�Z � ��Q�I�I�I�E�� � �?�0�!�,�$�0 ��@�O�^�S�[�O�����������      � ��?��������                                                                                                 �  g{g � ������������� � � ��8���8��� � ��� � � � � � ��8�\�m�~�}�{�&|�A�!�� � � ���8��<�x��D?Ŀa������8��� � �                                                                                                                                                                                                �W�Z�_�o�w�8�� H�E�@�`�p�x�� �� �&�6� ��U�?�@_�Y�I�� � �@�?�?  � � � � � � ����������������                                                                                                 � ��8���8��� � ��� � � � � � � �  g{g � ������������� ����?����?=���<� � � ��� �� ��`�k������Ө�Iv ���!�"�$�@�����B�N�f�:e�>�w�` 1  	      � �{�w�b�F�Q�Q�R         D�|���}��|�9��� � �           O����������L�}�� � � � � � �    �� �m�j�m�v�j�j           ���0Oϰ�@���     0 @ �     � ��@�@�@�@�@�@    ` ` ` ` ` �  �  � � � � �   � �           �?��y��=�}�u��        
 z ?�_��s�y��l�l�d        p      ��?���_��?�?         � ��x�s�g�o�o�o           ����������������� � � � � � � � ���������������� � � � � � � � � ���|�{�w��             � � � � � � �� � � � � � � � � �M�!�A��6�6�U�A  @  * I I *  ���k��x�i��2�V      `      �A�I�+�^�c�?�@�          @ ?   �X_���?����           �   �Y�Y�Y�Y�Y�Z�Z�T        ��3�'�/�/�/Я�                �@�@�@�@�@�@�_�@` o o o o o   � � � � � �  �    � � � � � � � ���������������
   ; ? ? ? ? �`�`�f�f�F�c�8�     /     �_�_�O��?���   o      �c�`�p�x����              �^�F�w�u�z���             ����������������� � � � � � � � ��������                 � ��g�N�]�{�w�n                � �o�i�i����  ` f ` ` ` ` ` � �o�n�n����  ` a ` ` ` ` ` � � � � � � � �          �  �����  � � � � � � � �K�W�\�B�[�]�J�l         Wh��Oϐp����p� @ 0  � �  � �� �7�0�0�>�?�    0 0 > > ?    �� 	�	���  �� �        �   � �{�t�d�D�S�P�X         � �@�_�_�_�@��@  ?       ?                             ��������                �oP� ���W�k�k�c             ����������������                ���?��� � � �                 �����������?��                ��	�o�i�o�v�I�O` f ` ` ` p y O ���o�n�o��`�` a ` ` ` � � � � � � �����    x p `     ����������� � � �        �g�s�y�|�~�7��           H p   ��5��������              �;�a�@��1�`�0�   > ` N    ����������          � � �V�C�b�p�x���             �^�\�Y�S�G�@��               ? ?   � �                 ���?�?������                �g�k�l�w�h�_��             � � � � � � � �                 � ?                           � � � � � ?                   ��������                ���6�����v�����                ��/������         � � ��       o � � � � ��������� � � � � � � � 8�����x�<���              ` �l� � �w�������               ��������          ??� � � � � � � �   @???  ��� � � � � � �   ���C�y�|�~߿���� ;    � � � ���������Ii�ͻ� � � � F �     �(�W��� �@`�>� ' o `  ?    �#U�t�0Po���  � p � � �     À�x�~��b��� ?   x � � � � �@� � ��  �/��             ���� �� � �              j��� �� �� �          � �   �����o�w�8�?       @ @ �p�{�;� �  � � �p { ;           ��������� � � � � � � � ����������r :  � � �  : _�U�U��*����8                �:�u�7���55    � �     � � ���@�?���`��_�? ?             � �������@�           N � ����ֵŦäۼää� � � � � � � � �[�kֹeھG���3          � � �
6�� ;����p�          �2���6�,��51 � 2 � �  ' � ������c � ���< > ~ � � � � � *ށu+��Ww߯� � ` � � � �     ���/�[�3�}�� p ` @          �� �� 2��m�-� �       M       ��������           � � �������`� �   � � � e  ����� � ���           7 7 � � ��=�9�0� �      = 9 0 & / U��*�
?���|��              � ���� ��� � � � �    n ` ~ � �?�?�?�?�?�?�?         ?�� ������ �  � � � Y    ääääۼääѲ� � � � � � � � �d����|� � �      � � � � � �  ��  �� ���               ���:���7�	        
 � n�gjwvwrwr;9 � � � � � � � ��/h/hH��G���� � � � 0 0 p ` � ���~�A��~�A    <     <     ���<�{�~�}�{�w          �  ������  �����    � �     � � ����������������� � � � � � � �                                                                 ��K�x�{�x�x�0� x 0             ��������               ��~�@���	��<              �o� ����� �m�m         @     ȹļ������������ � � � � � � � � `�?@������  ? � �         � ������ �   � ( ( ( �     � ������ �   �    �   ��|}xy�y`a;��� � � � � �   � ��� ���� �   �        �  � �`�`���� �p  ` o g s x   �p���1����  ~ ~  7 ; ; ; OH��_��	>?�     0 � � � � � �8�g������k�  8 p        ��������p p p p p p p p |������� ������|    �    w��w�w�w�7� � � � � � � � p ? � � � � ����� �     ?   ? � � � � � � � � � � � � � �  � � �B���X��?����              � �P�i�>��/�w�v             �w�v�v�v�w�w�v�v           ������o�`�@��       O �   � � � �    ��� ?� �     � ?   � �E�U�Q�Y�M�E�U�Q: * . & 2 : * . � ��Q�Y�M�E�U�Q    . & 2 : * . m��?�O�o�q�~�w�w             � ߿��7�������{             � ����އ��������    > > <     �΋�OH��H��	��0 p �   0 � p � � � �  � � � �  � � �         � � �    � � ��   � � �         ��������p p p p p p p p � � � � ����� �       ? � � � � � � � � � � � � � � � � ����������������� � � � � � � � �w�w�w�v�v�v�o�o             �o�o�k�m�W�'��            � ��hw�  ��� �     �   �       �����P�V�D�E�Q�U? 0 / ) ; : . * �T�V�@�F�@��� + ) ? 9 ?         ss��  ����� � � � 1 �       �!�s�y�|�|�?��                c� � ��   �� ��        �       �2��6M�����    0 �       ��v��}�n��� �         �     ���������������� � � � � � �  c�3��{vvvvv   � � � � �  ���?p�?� ����      � � �     ���������������� � � � � � �  ����7�o?���� � � � � � �  ����������������� � � � � � � �                                                                 �x���p�� �@�~� x � p          �~�~�~�~�~�~�~�~                ����s缳߹o�w�wh � s � � o w w ���<{Ͻ��{���s�� < � � { � � � 8�x�����������x�   @ � � � @   `�������������x�          � @   ��~�>����w��� � � � � � � ~ � � � ��� � �  � ? � � 8  � � � �f~�� � v�� �   w �   � �   �J��U����;o���~k � � � � � � � ��x�?�<�8�0�0��             ����x�0��8�x�              ������������       @ �   ����������P             ������7��8���� � � � � � � � ���~������� � � � � � � � ?�a�� �����z�|� � � � � � � � ��{^�?�a������� � � � � � � � � �$f�>�\�~�>c� f � � � � � � �9��n�7�7�g��8?   � �   ? ����������?        ��@�?��O�9���  ?       @   ��@��?�?�?�?�>  ?       �>�� �@���~�   ?       � � ��$�F�H��� � � � ~ ~ ~ ~ ���T�j��� � ~ ~ ~ ~ �    � ���D|������ �D� 8 � | | � � � �_��|���|��_�_' ?  �  ? '   ��������~ ~ ~ ~ ~ ~ ~   �  AAAA���  � � � � � �   � � � �@�>�`�p�|~ ~ ~ >      � ����	�	��   � � � � � �   �� � �
�N�_���       @     � �� �G�O�Z�\�W� � x ` @ A A @ �S�Q�P�X�L� �� D F A @ ` p � � � �?�s�g�F�^�}�s         � �g�g�g�g�g�g�g� � � � � � � � � �������������� � � � � � � � �`�`�`�`�`�p�� � � � � � � � � �������� � � � �  � � � � ���`�o�o�o�o� � � � � � � � � �������������� � � � � � � � �o�o�o�o�`��� � � � � � � � � �������������� � � � � � � � � � �� �@�@�G�O�_� �  p ` @ @ @ �_�[�]�_�O� �� @ @ @ @ ` p � �  �W��0�8��L�o�  ( D    @     ���-��(��   $ �          l�T�$�O��s�g� �   @              � $C���� �        � C $   H���� �@� �P�  @         @                       ���� �'�/�/�/�/�? ` @ @ @ @ @ @ � �U�U����U�U  I A A A A I A � � � � � � � �    @ @ @ @ _ _ ��������~               �  � � � � � ���                �?� � � �  ���� � � � � �    皽 @�@��?����;  B "    w                             ? ?                                                                                                                                                     � �������                � �~�}�{��?�\�l       ?   � � � � � � � �                 /��@�?��O�9���@ ` ?       @   �]�A�|��[�@�� A A   C @    � � � �B�_�@�� _ _  B C @    ��������                    ????????????� � � � � � � � �@� �o�\���M�f?      F F "  ���@�@������:t     " B    ���ke��
�
c��   � h d   ������ � �           ?     � � � �  �  � �           �     �d�C��b� p�7��  8 `        �����
��� �    � �     � � � � � � � �       � � � � � ��� � ����        � � � � � � � �            � � � � � � � �    � � � � �     8 _��8   ?h7�|�x  � p`Lp���a��   � ���:����x                         	           �          �0        ` � � `�        ` �`�`��                       �               �                                         � @�@           ������  ~      ~      ~      ~      <   <          <   <       ,Z�8�4�d�l  4<f~��������� � � � � � � �  ���������  ����� ���������������< B<B<R,B<B<B<< <<B~B~J~Z~B~B~<<   $< B<�~�<�B  <<<<B~�������0~"/       �p] , 
       �� � ֔���     �@�@�@j  �     
  	   ,�<�� |��� @�� �����0|0<�� � �         ` � � `�        ` �`�`��0             ?             ��|x00     ��D|Hx00                @ @ @�@��       ����������           
 
 8 8       



8888                         �t�d�h�X~ <    ��������B~$<  � � � ����� ���x�p�`� � ������������ ��������� � � f�f�D�^�~�~~ ~~����������~~�~�f�f�~B<<     ��������B~<<           ??       	  ( 2       � ��������      �   P P                       
         p �@�@�         p h h �   f �f�~�f�f�~r<  ff����������~~      ` �@�`�pz8      ``�����F~           	                � ����        ������                    ff�߫���bb44   f �T�>�~<     ( |(|8l8(((  ((T|T|T|888888(((((D88  8888888888||(8    
 
6    

*> <8     $<'?          �                �        8 (4
 8 8 <     ?/ * 0 $   ; ? /   ���@h h ��8��� ( � � � T � h � ".5
&>   ; ? ; 9 9   ��쐖hV��44�� � d t � � > � � � 44<2<2< <<<<<<>><<>><<99z8�p�`�@`   '?'?F~������``           ��� � � �       x���������           ~ ~          ~~~~    ++uq��~~   ?
<� ~     8 8088       88G??G88          �  ��           ������    (((((      8888888888         ���       ������    � � � l6 � � � | >       � �@�03      � � � ?              ����p�8�����    ����������������������������������������������������������������������                ?      � ��0 8��       � �������        ; <     ??    �   � � � <     ���`� �h���   $J4^(<      <4~(~<       8 ,         8<     �������� � �0�8������  � � � � � ��� � � � � � � �������������������������������������������������������������    �  ~ <     x�2$~<   @@         @       @"  	  @@""  		   d����  dd����  ����������������������������������������������������������. . <1  ???? t t <���  p � ������p�@����� �??>?    ??	??   ��|����@� �   �� ���8����� �  8 D8�|��b~,<  88||��b�,~<    6~ Z4d88      >~,~| 8  ���������������� � �?�?�?�?�?�?��������������������������������������������������������������������������� G�B�p�pp     G � � � p     9l8�x�xN0;    9 | � � ~ ? < v4< 4r<�bv4< <<J~<<,<~~��J~<< x � �@X v�b�bhx����xxn~����  ~ �b�v~ <44  ~~����~~$<,<,< 8 L0((((((8t|8888888888           0 � � ���@��    00����`�����    ` � 耰@��(04| ``��x�����88<|           


   ? > ?  ?    !?.>!?!?  .      .   ..QUUUQ..  f �f�~�f�f�~r<  ff����������~~    ? ?       ????    � � � � � �     ������������         
9      &?  ` � � �@���|   ` �@̰�H�����8 l(�t�d�Pw(6 88T|������Y>>�z�d�@l +% ������t|5???~ v<�B�~�B�f~<< ~~~~��������B~<<(l��T�T��   88||����������  2f8�x�p�rq9? >>x~������??48:�u	��� <<>'�w����??t<r:9 2?8?||~~??� |
��8���� $�|��������   > > ?      *>*>!?
   ? ? ? ? ?    !?-?!?-?!?#� _@_@���� #�  @�@�44<2<2< <<<<<<>><<>><<                                                                <;8   #?$?'?  ,��80�����   ��$������0���       Tl         l                   
          0 0 ` `                                              ` X,7                7��|��M�        < � �   >!>!A^cLw    ! ! A c w   ppȸ|�|ľ�r��  p � � � � �      
              	  ��p � �     0   0 �       0   -3>!~A]b     3 ! A b   ��<,&:������   � , : � � �    /<8/p/p        0 0 88L|�Φ���||88  8 | � � � | 8          CC�G        C         ���`�D�         � � �    @ (         @ (           � | 8 | D    � | 8 | D   ��Bf<Z$<$<<ZBf��� B  < <  B �        @   � �      @   � � '.        �|k���K��� � t � � � t �     $?%>? :%  ? >    %     �<��&ڄ���    <   � � �      3! !       @                � � @ � � @    � @   � @       !?    ?          oi��T|((66hX00 i � | ( 6 X 0     (8           8            4,,<         , <      ?>?*u08    5      @�x�<�<�L��8 �� ` ( 8 H       oG�!v&     e "      �  ����x�        � p   <~.       .         �@�ހL�``� `    � �   @                      � �    �                    �� D (  ( D��  � D (   ( D � (8Xl��h| 8    8 h � x         ;;|O��ot_n_n  ; O � � t n n  00L|�~����>J40 L � � � � J 4     	 "3             @ � � `������        � � � �   ``P`(1 �  ` ` 1    �  ( @�����p��p (  � � � | 0 ����  "DGP�@� �   D  C � @   (T` 4�T�    ( ` 4 �    	898          �0�p��\hܨ|@� �  `  X � h �      ?7       	        8(|���<�| �    8 d  8 X    � `Xx$<*6
� ` x < 6              ��@��`          � � `     DD (  (DD      D (   ( D       ��       �    WnyF?0P����G88n F 0 P � � G 8  � ` P(
  � ` P (  
                     �����p�� �     � � � �         �S�@o+\1~? � S � n X <  �  �8�ز���P@�� �8 � � �      � ` 8         8       
��  @P`     �   @ `      @@`0   pS pĠ  @ `     P 0 �      @��@A�E��    @ � A B  �   `1>� <3     >   3      �<����C���px  < �  C  � x     ���x�ZfZf-3    � x � f f 3 �p��Tl*6*6*6p � l 6 6 6   tl��h���p`��� l � �  p � �      (  (          (   (       31=<MDww?:~d Y  C �  �    .,91&&wu}i> , R  Y � � 1   ��<<fb[Y>.5 J 0 B � & Q <   *1JD      * 1 J D   �@ 0(    @ 0 (       p �Pd` "tF    P `    t F   � , b�p�x��       p x � �    JD��@@      D � @    lTF}*}m??' D | = ?       �6�l�$���X�d    l � � � H     ;=��:��<8���  = � � < � �   :(8*0
�J�n\d    ( * 
 J n d ~D�Ըƒ�:�ZfD|88D � � � � f | 8 &0P0 @ �  &   0 @ �   ""uW,?+478Op/0  " W ? 4 8 p 0  (�>�|�e 8 ( � � � e  8 ((@p��h�b�0�	�( P � h &    p����^�K� `o 0 � � N G # h 8px �P��\o
W�0 p ` p 0 L F # @l38  @ l 3 8      
n4��,�X0���   n � , X � �   "Ca(001   C a 0 1      d�D��X0���    D  X � �        @                             >   }       > 9 6 5     8 | � � �`��      8 | � l �     8 4         ,                $ t               � x �0� g9'     X � � `           '#        & #     � @ � �`�0�p    � � � � � � ! x���Nsb}=  � � s } =      |@pLðB���    @ L � � � � ? `?����x�x�x? ` � � � � � �  !

�         L � � ,��<��v�    � *  2 � �  !

�         @ � � 8��2��v�    � 0  < � � '+~&�O�5�)^I� # Z �  V N � @�0��=4΀��:�� 0  � � 2 � � <>                <�|���� � � �   ( X � ` � �       .Rd �``    2 n \ � `  v?>,vZ�~�<f <$   4 f B $   �  �0� e9'     P � � e     !!!	   ! ! !   	    ��H������ ��   � � � �    �   
   x        x   ��� "@8`� � � �   8 `        ?�         �     J7-           5          ���0���@j ,  � � � � � ^ <  J7-           5          ���0���@j ,  � � � � � ^ <  	��٥ߒowF� � � / ' G   �>�߷�j�����| � � � � �  x   ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �                                     � �             �            P l{4          p | w          
6�,          > �      337       ? ? ?     � ��~D;����    � 4 � � g     
              � �`��,�p_��  � � v r � � �    >     ? O K X   � ��0�<���� ��  � � � � � � : ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �  ��������������� � � � � � �                  � ����x|8|8|   � � � � | | |   �c�h�	��n} � � � � �    =���� �l�r�|| � ? ?  � � � | 7?   ? ?        � ����0p�� 0 � m " b � � � 0 3?/&    ? ? 3 :  ���l���`� �     � � � � � �     ��A�dw	> � � � z /    ���^ |0 � � } � � � � � �    /7s      ; , O   � ��0�8�����0  � � � � � 4 �    ?7       # *   � `�x������8�p  � � � � � � r           P l�t          p | �          
6�.          > �           0 H0w          0 x           
�           �             8 '            8 ?            4�0           < �             8 '            8 ?            4�0           < �  0g8�p�`� �                � ��������             �8�?�8�;�;�;��            �4�����������       � � � �   ���`0? � � � H 6    �y�����p��� � � 	  l � 0 � 3?77]8 - 8 / , z '   � � � | ���p��� � � � � d � 0 � �c�(�I�L}- � � � �  ?   =��m��4�x�x�pp � ? ? { � � � p �s�@�{7< � � � O ?    <���<
�4����� � > � � � � � � K5V)v	[$j4; G O o   ?   ��x�x��z\�0�� � � � � � � � � M3Y'w7/	 G O  ; 9    � ���t��ĸ�0�� � � � � � � � � �9�
�e�b�a�p�8�8              ��y��C�`^�*ՙf�7               W/X'_ [$K4c0                 ���������                <6>}"    ? ? ? ~ � ��� �0��(�8�� � � x < l | >  8 ; lE:L7, ( + _ _ ~  ?     � r̹n�.�v�    � �  ?  �  :~      ?  � @��@� ��(�|�.؀ � � � � � � �    /s,]n)     1 ]  W ~ �B�������~��~�~ � � � � � � �      /3}"       1 = _   ~ �B�������~��  ~ � � � � � �     � ������0�D    � � � � � �       /3        1 =   ~ �B�������~��  ~ � � � � � �        , < $ 4        4 < < ,         ` � ��        ` � � �            ��(           � < ^#! 7   { y >    z������X0�� � � � � | � p � ??_ 0w(: ? ? s O _ ?   .�����,�p|���� � � � � | � � � _/.~=<    ?     ���t~�<����0�@� � � � � � � � � 17    K ;        $����ý�<~�<�� � � � � � ~ < � ^o)?  g W +      ~�$�����=g��X� � � � � �  � � z�����@Ȱ� �   � � � � � � �   =o-/';: / S 3 ;  ' &  ~�$����ý�<�� � � � � � �  � 444 $        , , , <        ?_%L0~ ?  ? ~  s 2    <�������@� 0�� � � > ~ � � 0 �         ` � ��        ` � � �            ��(           � <         @ � ��         @ � � �           p �0�P          p � x      ={$_O	      # ] g w         ~ �~��<�        ~ � � �        ={$_        # ] g           ~ �~��          ~ � �       0 X �@�$�      0 h � � � 8 < z4][O /	  < N k m  7        p �p�~?���      p � � � �  8  T T |                        D � D                          < f$�B� �       < Z � � �  8 llllll ( T T T T T T     ?  �? ?       ? @ � @ ?   ?_%L0~ ?    ? ~  s 2     <�������@��p� � � > ~ � � � � ���~}3{A>> � � �   { A > x��h�X~������   � � � � � � �   /	    7         �����<~��~�<<�� � � � � � � < � O	/	    w 7        <������;{�ƽ�? � � � � � � � ? ����@P��  �� � � � � � �   � �                    ���?�α�= � � � � �    8 (((((((8 ( ( ( ( ( ( (       � ��           � � �     �$��Z $      � � � f <      | T(D8(| D8( D l | 8 | D (      � �d�6�d�       � z 9 z �        /?^#_1      7 7  {      (�0��z���     8 � � � �        /        7          (�0��x�       8 � � �    /    7        (�0��p�����   8 � � � � �  / 7 ?      ?     � ���������    � � � � � �      =6        ?      � � � ����m8    � � � �  �      =6        ?      � �`�0����}8    � � � �  �    //7    >   ? /       � p�8��(��      � � � � �   ??~7     ? ; w � ��� `���� ���� � � � � � � � �m�C��K     � � � � O 
    ������u@� p     � � � � � P     ?''36 ; = ? ? ?    �����̸l8�0x0 � � � � � � x 0 73   ? ?        ��̸�p�p�0p     � � � � � p     ;7	 7 ?       �0��x��������� � � � � � � � � '�o�~     w � �        �<�|�������     � � � � � �     '�o�~       w � �         �<�~���88       � � � � 8       .?	?	?   ? ; 9 -      t������������   � � � � � � �   |??      ?        �x������ݸ�t`� � � � � � � � �                                                                   ??~7     ? ; w � ��� `���� ���� � � � � � � �   7'      ; 9   � � ��:�~���  � � � � � � �  .'/    ? ? ?  � ��p�8�t����xx�� � � � � � � �  ?2�c�g|?~  ?  � �       � � @�@�@��     � � � � � �  ?13>?   ? y s ? ?   � ���  � � �@�  � � � � � � �    <x���    3 W � � �   � ��|0�O    � 0 � 
 � � �       ` �`�`�@      ` � � �         ���         � �                                                                 |??      ?        �x�|�����8�t`� � � � � � � � � /.   = ?       ��t���� p@� � � � � � � � � ` � 7      ?   x�p���8�p�� ��� � � � � � � � � O~? _  O  w '   � ����m����   � � � � � �    ??'> /  ' ? ;    � |8n<�t��5���� � | ~ � � � � � �w5:;  � J / $     �T �����  � Z � d   �  n=n;>8       ? 8       v�v�<����       � � < � �       �m�a�]�>����]e�A��>����]����k��x�i��6�V������r�`��T��`�s�_�o�?e>	w,`�3�W�O�'�	?$    ? ??=;?     ??????@ � x > =   	 @@��Xx&>#?    � �0�:�y��  ����������  c �  ?    �?? � �f�B�f�<� � �  �f�J�f������� �  ( ( h h h �   880x0x0xp�  4 : z z } �  <><~<~>~�  8??????  88????????????      ����������      ����������                                ����            ����1111! !//????? ? ? ?L L L L � ���xt8���������� � ����I�I�+�^�c��� I�I�*�\�@��� ��X_���?����� P�B�
������� �    ���  ���        �� �����     ??� ??�? {???G??����?�����o��y�����������������      ? � >          ??�?       � ~<= � �        ������� �� � ����� � p�`�P�P�P�P�`�p�� ������� p�n�Z�P�T�Z�n�p�????1     ????????1?     �����������<� ����������<��               �����������     ���������� �    /�_� �@  ?    ��?� �8� � ~ ��� �� ������������� ������������������������������<<B~�ý��[g~Z$$<<~~������gZ~$$�$�$�$�$�$�$�$�$Z�Z�Z�Z�Z�Z�Z�Z�,,vF����nn<< <~\�8�~ <  204z   ???E� ��8 <0< �� � �����������B�ǂ�B@?@?�?����?��B�" ������A�B��������A�B�D�H� ������� 8?8???????????????� �����<����x�8����������������                       ������          ������               ? �;����������  ??������� �?�?�?�?��!^�� ���@�H�^�!� � �� � ���䅄{�  �������z��� �������������������������������$�$�$�$�<�~ < Z�Z�Z�Z�B�f�<~ <8 D8�|��f~,<  88||��f�,~< 4,4,4,4,4,4,4,4,,<,<,<,<,<,<,<,<��Lo0 ~?  ����{~S/?����� ~�� x�� �����~������������@?@?@?�_������ "B������������A�@���� ��D�B�A�@�?=???> ????????????�8�x�x�x�xl���� ����������������              �����������00   ����������0� 0  ???x8`  k6k6 ? ?@G_ww������
����������@ @ @            @ @ @                                                                                                      P(V�R([([(\( �<  �,�, � �  q(   �(�(�$�$�h�h      T(�<X(�,�,](�$�$�$ �$�$ �$�$ �$ �$�$�$           T(�<X(�,�,](                          T(N<Y([�[�\�                 %%       T(^<Th                    %%       P�V(P�                                                                8888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888       8888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �<�<n$o$�<�<�<�<�<�<�<�<�<�<�<�<�<�<�| �<�<�<�<�<�<�<�<�<�|  �<�<�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�| �<�$�$�$�,�,�$�$�$�|  �<�<�$� � �$�,�,�$� � �$� � �$� � �$�| �<�$�$�$�,�,�$�$�$�|  �<�$�$� � �$�,�,�$� � �$� � �$� � �$�| �<�$�$�$�$�$�$�$�$�|  �<�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�| �<p%q%r%s%t%u%v%w%�|  �<�$�$� � �$� � �$� � �$� � �$� � �$�| ��������������������  �<�$�$� � �$� � �$� � �$� � �$� � �$�| �(�(�(�(�(�(�(�(�(�h  �<�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�| �(!%"%#%$%?%�$�$�$�h  �<�$�$�$�$�$� � �$� � �$� � �$� � �$�| �(�$�$�$�$�$�$�$�$�h  �<�$�$�$�$�$� � �$� � �$� � �$� � �$�| �(�$�$�$;1<1�$�$�$�h  �<�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�| �(�$�$�$=1>1�$�$�$�h  �<�$�$� � �$� � �$� � �$� � �$� � �$�| �(�$�$�$�$�$�$�$�$�h  �<�$�$� � �$� � �$� � �$� � �$� � �$�| �(�$;1<1�$�$;1<1�$�h  �<�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�| �(�$=1>1�$�$=1>1�$�h  �������������������������������������� ��������������������                                  �$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�d �(�(�(�(�(�(�(�(�(�h  �$��$�,�,�,�,�,�,�,�,�,�,�,�,�,�,�,�d �(y$z${$|$�$�$�$�$�h  �$�$�$[-X-U-c-'-�,a-T-P-S-�,c-P-[-Z-�d �(d,�,�$�,�l�$h<h|�h  �$�$�$�,�,.,�,�,�$�$�$�$�$�$�$�$�$�$�d �(u,%=�$�,�l�$x<x|�h  �$�$�$_-d-[-[-�,�$�$�$�$�$�$�$�$�$�$�d �(�(�(�(�(�(�(�(�(�h  �$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�$�d �(i$j$k$l$m$n$o$�$�h  �$�$�$� � �$�$� � �$�$� � �$�$� � �$�d �(�(�(�$�$�$�$�$�$�h  �$�$�$� � �$�$� � �$�$� � �$�$� � �$�d �(�(�(�$�$�$�$�$�$�h  �������������������������������������� ��������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���u��u�u����������������8�������{���K�{�������{���������n��������������������n���������n���������������������������,���������t�5�T�e�u�t����� ���{�����;����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;��s����������������������s������#����������������������������������������������������������������������������������������������������������������������?���������������������������������??��������������������������������������������������#�c��c���������������������������Ϸ�����������������������s�y�9�1�������������������������������������������W���]�=�����������������}�����������������������������������O�w��������������������a�����������������������������������������������1�-�����g�������������������������~� � � �����~� � � � � �~� � � � � � � ����������������      ��E�J�w�n�^�����      ����#�&������g���k�������								������������������ � � ���      ��������������������������������������?{�g�_���          �  ���          � `� ������������������ � � � � � � � �������������~� ��������������������������������������������������?�_��y��/��������������������������ߧ��?������������Ɛ���?��?�����;����������������������������������������m���������{�H�k�����������������������������?�?���������D�m�l�m�l�������]���U���]���������������������?!?-?-A���``����������������o��������?�?����������������������������������������������Ǹ���?��?�����������������������������������������Z�Z�Z�����������������������������Q���������������������ż���?��?���a�9�                ��������������������+����}���{�����������������������������������������������������������������  88Gx_'?>"�����          	�� �࠰P�P�� ������������������     ???        ��h�-��M�m�������������ƻ�������7�w��w����??���    ���           ?7"n"n|xx  8|xx  ?2>?~ll  ?2><2>"n|xx  7?2~f~<88  ><2>|xx  <~"n|xx  ?!gBN800  ??2~"n|xx  ?7>2>|xx�������������������}��G�I�I�S�S     |      �����������������#������Ͽ���?����������������   66I>A>A"   66kUk]c*6   66>>>    *""     �������������������������  88G_x?'">1/gYϵۭ�����������        ����������������"f"f"f"f"f
~~~  �w��w�D�A���  �������������������������������������������������������������������ߣ�%�w�ß���������������������m�s��O���7������������������������?�o���������������������?s�9ϟg�3�����������������������������������������������������?�?������������������������?��������������ݣ�w�oן��������������������������������o������������������������������������������������������������������A=�c�����������������������������������tLtLtLtLtLtLtLtL�������������������������������������?�������������������������/�/��?�������������������?�ܿ޿����������������������������������������?������������������������������������������������������������������������������������������������������������W������������������������������o�o�����������������������������1�y�y�a��������������������;g�{���M�U���������������������?�����������������������_���'������������������������?��_������������������������?���?���������������������������?��������������������������w��������������������������s��������������������ߺ�������ÿ�?������������� ���������������������� � �����  ??DoPrOsm~J|D  ��� �  ���    ��������������������������O���  ���������������� �  ���������  �� �� ���&���?0wHxGׯ���������������������������������������������������������������׈��ܫ������ �  � �� � �� "B=�?�?��� � �q�Q�J�U�[�� � ��0X W T#W  � ��4�U��� ������?F8�p�8�D��B�$<D|��d|$<$<$<<<B~��������io">">">R~R~~~�������������">$<D|Hx����~~����y	<<B~������������~~������������������������������������3 8h`�� � _��
Q�Q���?�pp P W T#T#�# �q �U�U�w���� � �������r�����������    $<$<$<$<$<$<$<">$<HxHx������~~R~��������r~��io	io����B~<<������������B~<<<<B~����������B~||������������������������``��������������||������������������Z���R���Z�������9�������6��������������������������������a��������������A���������������a���������������A���������������C��������������������������������������o���{��������������������������������������������������������������������������o�o��������        {{J{J{J{        ��	�	�y�����U���o�l�������F���l�m�m�������n���.�����������?���?���?�����        HHI�����������s���        ��$�$����������������������o���{�����������������������������������������G�������������������������������w����������J{J{J{J{NBBy���t�z�
�
��������������������?�?����?�?������������������?�?�������������������C���I������)�(�(�����d�d�����!�!������������������������'����������������߸ǿ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������}�9�U�m�}�}�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������j���������q���������������������������������������_���_������z��z�z����������������������������������������k��������� ���o�����/�������m�m�����^�����������������������{��s�{���������}��������������������������������c�o����������o�o��o�o������������u�u�����c�����c�����������j�j�j�j�����������������c���        y �0�I�A        � :��%�%        � �F�I�I        } �(�1�!        � 0�� �          


        � �F�I�I         ���   � [�[�[�  � h�h�h�h�h�h�  p P P \ W(K4[$        � �`h�h�        w U"U"]"        { �1�I�I        � �Hu��        � C�B�B�   

�;��$�$        � �am�m�        � y��I�	          � � �                 �1�	�I�I�0y     ���%�%9��     �O�H�I�Iy��     � � �!�!� q     0�� � �&9�� 



	     �O�H�I�Iy��     �����     [�[�[�[��D�     h�h�h�h�h��     [$[$[$K4W(<     �x�h�h��`�     k**6     �y�A�I�I�1{     ������ ����      ���$�$;��     n�o�m�m��a�     p��H�I�Iy��     � � � � �                         p P P � �x�!R!        � 0�� �   x �0�H�H�@�A�0        � :��&�$        � �m�m�  p P P � �y�!R!        � �#�$�         � �g�m�   �V�V�v�  � � � � � � �                                                                                                                                                                                 R!R!R!^!g=     � � � � 0��     u�	�I�I�0y     ��$�$�d[��     o�o�m�m�s��     R!R!R!^!g=     �#�$�$�e]��     i�h�h�h�h��   �Q�Q�P�!R!� 0�� � � � � � �                                                                                                                                                                                       � �@�@�@�@�A�A   �8��"�"< $$4�{��        � 0�� �   � �@�@�@�P�i�I        � 0�� �         y �0�I�H        � :��&�$        � ��$[$  x �0�@�@�B�B�   		�	�I�I�I  � � � � � � �                                                                                                                                                 �A�A�A�A�x�     ���"�"6��       �C��     0�� � � 0��     �I�I�I�i�Py     �� � � 0��     �@�A�I�I�0y     ��$�$�dZ��     C<^ Z$Z$f<     �B�B�B�B�A�     �I�I�H6ɶI�     � � � � � �                                                                                                                                                                                       ��V     �    ��    �i�    ��9    � =C     8�   �    c��!s>9WN��c��!s>9WN�  �k-�R�w2%��%�c�-�+�  c����M}{�c��	�+�  c�0*���$�c�S)Bc+�  ���5�s)5��Y�c��	�R�s  c��&)}���c�  ��  �=;�fR�B)&�Yc��!s>9WN�  ���J�?�  �y��9��f�E  �Ii�b�o�QO~  �Z�U�v��*�  ����6��A%  �������  ��1��6�V~�e  ��IS;�_7  �~#u�6�q`  ��'-^��z�d  ��2� >&��V�9  �k-�)�/%�w�R  �~#��6��x�YG6h;J
�\*qz� �`    � �8    x �8    � �  � � � �   � �  � �  � � � �4   0 �   8 �   � �    � �    � �8    � �    � � � � h � � �  m �   � ��    ��  ���  P a�    Q�  G �   [ �   G �    J �  ] �  e �    b �   Z �  � �l   � �    � �    � �    v �l   � �    } �    x �    s �    w �l   q �l   q �l   n �l   � �F  v �    v �"  K �  [ �  k �  { �  K �  [ �  ��   0�    v �    v �   ��    ��    ��   { �   (�7   0�8   v �l    ~ �l   | �   | �"  8 �8  @ �7 ( �7   0 �8   8 �8   @ �7  ( �7  0 �8  8 �8  @ �7 � �D  � �D  � �g  � �f  � �}   � �m   � �~   � �n   � �n   T �B U �B b �  x �    x �"  e �    e �"  r �&  I �M  < �l   ; �l   ��    ���   k 7    l >   ��     j�     j�    t ;   ��    ��    m Gl    u Gl   l 5   l ?"  c �   c �"  x �    x �    � �,   � �  � �   � �   x �l   � �  � �   � �    �         �                      � U_�N�                 J   �Ҳ��������U�  N���     �   �  �� �  p�           
.-
.,"                                                                                                     13                                                                                                                                                                                                                �I�I_�                                                0�`�$�@0�`���
��
���
�
 � ��	 ����������	�ܦؐ�٧�?ٹڷ�Y���R�                                                                                   � �                                                                  � � � � � � � ��@  @�       �K�$ K�K�K : $ <     
                        
  
 
 )  $ &  0 + -U   ������ #   7 & - - 7 < �!�$�!#&�!�!j$I                 ` $   $   p�   � �              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �Ͻ� ]������ � =��� =���?"�H�`�?�	�?�	�<�]?�	���� ��� �S��� �
���iML��L���� ��]��� ���E�F�D\\�kk�� ��m�8�`�C�C�1?E?m�?�?�?��?�??��?�iML�����\��L�S��`�Q�Q�?�
� ?�_D��� �G�1�?�==G��_D��� �� u� ���� ���� � o� o�ʐ?f���Ȱ��$G���(`�P`���a���`��\� |ՠ� ԰� ����	G^	GE��Ԡ���ԡ���
�a����a��`�a?�?�� ���4�	�����z�M�� ��]��������-�����ݍ z�+�/K|=������ ���� ��m�!��z��!����z�}�\��?�	��-�G$���� �� o� �,?�	� �<?�	���\?�	?�� ����������ò�Z��� �[��Y?��\_ ����Y���p�Y_ ������Y� ��_ oh��h��h���h���h��
/$���_�H�F � � Go� �@:@-�@:@��o`� �����]��������@��H�F o���G����
?��Ձ��Հ��Ա��KG���Z�h�T�P�B�_��Y� So� �_c
������_y
��]n�?�
�%��_�
h��h��� �/�B�B?�
�B���@/�����0 ��� �G�1�
��� ?f� ԀԐԑ��p==G��� �^�G�D�1�z�p�l?\����?������0�0�1�1/�0 � ?\0-�(���=��(���=�?\h��?J/�����-�G$��?	� �p�������q/��?�?z==G�_t�T��VzRnT�T�R�h��dz`�`�fzbnh�h�`�j�b�Z��\zXnZ�Z�X��^� �G�1�??==G��o��+-�*-�\�����0�0��1�o�����`�_���`� �=�$G�:M}�\]� �(8 HH 	GI�/�GNI ��� �� =�������!��� o�Q(�1� �0oԑ-?\�P��1�?��@��Aoհ?\ա?\Ա��� ձoձ-� ��Ξ�D��o���	���� �Xo�Z?\�[��Y�Z?��\o� �Ro�T?\�U��S�T?��Vo�Po��o��?\��?\��o�/� Ր�Ձ?\Հ?\ՑoՀo�� � oԐ-?\� ���?����oՁo�@?\�A?\Ԁ�0�0�1�1�@�0�A�1o���J?\� �`?\� �b�Ho�h?\�i��a�h?��d?\�j��c�h?��fo�`�b�Ho?"?\�N?\��]���?�	=�`����Do�M�}�� �� dM�+(H��L`�L�L����� � �� ���H �l?�	�M�}?�	H���Ѝm_�	�_o?^o���o��_�
���D�0h��>�G$��?^n�/-?^?\ԡ?\Ԡ?\`�P��(Հ��a��m�?��p��qo�a��`�o�kH��� �-� ���D����of����.3EHLXy���[_u��� ��h       ���	� ���?����#����	G^�����/`����?[/����?f���	�0���?��G$^�F�1��0�}�\���y��x����`�x��!��QݐH���?�	�� ���3�o	G^��M�`�
�� ��/	�?�����o�q�e�q���p\���0�1�� ��0�0@��h��?h��)h��0m���@�/���#��
�1-�0�/��A-�@�/���-����/��G�\?�	���������/�$G���`���?�?����L��ްD� u����/@�  ����`��Ա��`��ՠ��H����h�(�/�ݍ ?F_l	����o����	����?N�1��0����
�A��@?0�?��?�������
�q��p?0�����ް��Q����`��_���?�m�Q��� �Q��z?�z�o��Q����`���H�����H��Y���������!o )4BQ^gnswz|}~       X����!++���43 ����,<MlL\=-\acNJHEIKF_�e	�	�
,��J���*Ver S1.20*��� ��� �� h���/ �� ��^� ��� �� ����/��^� ��� �� ��� �� �� ���1�� o�(?]�����̀����%��`����d�7��L���/3�(?]�����̀����%��`����d�	��L���/��/`�����&���L�\������������������ (���%����$J��J����J�M?�	o�����������\?�	?io�h����o� ����ՠ�ա� Հ����\?�	������o��ՠ�ա� Հ��@�\?�	��������?%����?%���o�0Ќo�����x��o�������?� �o\���p?�	���?�	�`��?�	���?�	_M��Ho��o��./:?`���(����(?ՠ�ա� Հ��������\?�	��]���пo��./:?2���(?ՠ�(����ա� Հ��������\?�	��]���пo���_������0��������}�\����� ������_�L��
�o�����ա�_|�����Ց�-��Ր�,_�����.��������}�\����� ������_�L��o�����ա�_�����Ց�-�Ր�,_�����.��������}�\����� ������_�L��o�����ա�_:����Ց�-�Ր�,_� ��ՠ�������%���������/��%���������/
��������D�?f��%��$J��J`���J�M?�	���������o��%����%��?i_:?i_|?i_�?���������,���հ�_�:,���\��� �,�0q��ֱ:,�,�0c]��%��.}����N���?�	� :,�,]����?�	}/5���?�	/(}���!�
�Q� � 
�
����� ?�� :,�,h��_Jh��gh��xh����_����?	��?�����հ������?v/�u�����\?�	���-Ց�,Ր��%����%��_:_|_�� :,�,���D�?	��?�� :,�,��ԡ� :,�,��Ԡ-� :,�,����D?�_�� :,�,�	�]���� >?�	=�n�� >���!� � _��`���?��a��`�� G_l	-�\� ?�	��L_�	                                  R&b&w&�&O(O(9'6'���b,>������$�    �b,>    
             &%&4&C&�%�%�%�%�%�%x$�&$$�$�#�#�#�#�#�#,#D#V#n####�"w%�"�"�"!�"�"�"D(R"�"?$3 ��� �G�� G�ogdCo��b$7�"�#5$            ?     >                =    ;  : 98    36                                                 ;            < N%J""�%�!="�!�!�!�!�!�!�!�$m!O!^!;!l$/!#!�%� 
%�� b� � K l'�'�& C �{@�&!���]�S�x�fs��� � v!�$�$�$�$              <;         8:       9         753     4      =>?             <;        :                  =>?�P�� �F�� �2�� ��� � �n� �$n� �
<�� �
F�� �
P�� � d�� 
��
}�� �}�� �� � �n�� �n�� �_� �P� �A� �-� �� � �<�� �F�� �A� �2� �-� � �x��� � <�� �� � � <�� �� � �
d�� �� � �
d�� �� � �(�(��4� � �(��� �(�(���
� � �(���
�� �x�� �� 
� ������f������f������f����x������f������f������f����p���<�����f������f������f����x������f������f������f����x��������f������f������f����x������f������f������f����p� �<�����f������f������f����x������f������f������f����x�  ��@�N�d�|�X�\�b�,�D�`�D�0N� �`2�� `�`*� `�`##� `�`(� `�`-� `�c2� `���02�� 0�0##� 0�0*� 0�32� 0���<�� �P� �d� �P� �d� �P� �d� �P� �<� �(� � �(��2��<��F��<��2��(���� �<�� �P� �d� 
� �0x��`� � �0x� �`� �  �0x��`� �(��(���
� � �(����
�� �P����0� � �P���� �
(����<����P����Z����P����<����(�������� �
d�� �d�� �d�� �d�� � �
d�� �� � �d�� �P�� �<�� �(�� � �(�� �2�� �<�� �F�� �P�� �Z�� �d�� �n�� � � d�� �0� $� �P��0� � �P�� �d���P�Z� � <��� ��� ���� �� }� �@<��@�� ���� �� }� �<�� �� � �x�� � �x�� �n�� �Z�� � �x�� �n�� �d�� �Z�� �P�� �F�� �<�� � �x� �Hx�� H�Hx� H�Hn� H�HZ� H�K(� H� �x�� �� 	�d�� �� 	�P�� �� 	�
��� �x�� �x� �x� �Hx� H�Hn� H�HF� H�K(� H� ������� � x�� 	��$� � d��$d� �(�2��
� �F�� �x� �x� 	� ��� �� �(� �� � �P�� �	x� � ���� �d�� �Z� �P� �F� �<� �2� �(� �� �� �
� �� � �2����<����(���� �2�� �<� � �<���$� � �<���$<� �P��������� �x���x���n���n���d���d���d���d����x���x���n���n���d��� �P�P�Z� �P�
�Z� �P�� �� �� � �$2�� "�� � �$2�� "�� � ��`� � ��`� �P�
�Z� ��� � �d�� �d�� � �P�P�$P� �F�2�� �P�� �� �� �� �� �F�� � �P�� �� � �x�� �� �� �� 
� ��� 	��<����2����(������������
���� �F�F�� � �Z�0� �x�� �� ��� �� ��� �� �� �� 	��d�� �d�� �� 	� �d�� �� 	� �0d� �Hd� �<�� � �
x�� 
�
� 
�
� � �<��<� �<�� �� � �2���Z���F������ �d� �x�� �	� � �(�� �<� �P� � �x�s�n�i�d�_�Z� �d�i�n�s�x� �x�s�n�i�d�_�Z� �d�i�n�s�x� �(�� �#� 	� �(�� �#� 	� �F�����`�<�����`� � �(�����`������`� �
P�� ��d�� � �(�� �� � �d�� � �x�� � � 2�� �0(� -� � x�2�s�(�U�-�U�-�U�#� ������ �<�� ��� �7� �
� �#� � �(����� �P�
�Z� �P�� �d���`� �d���`� �d���`� �0d�
����(��P�����0� �x���`� �d�� 	�Z�� �U� �_� �K� �U� �<� �F� �2� �<� �-� � �(�� �2�� �-� �� �� � �(� � 2����(��������
���� �(�� �2�� �#� �(� �� �� � �(�� �2�� �-� �(� �#� �� �� � �P�� � 	P�� � � P�� �P� � �P������ �P� �x� �
x�� ��2�� �-� �(� �#� �� �� � �F�� �x�� 	� �x�� �� � �x�� �� � �x�� �� 
� �`P �� `�c� `���` P�� `�`� `�c� `���`2 �� `�c� `���` 2�� `�`� `�c� `���`� � �� ���0 ��$ ���`�� `�3k� 0� ��� �� �� �� �� �`� `�c� `� �(�� �� �<�� �� �P�� �� �<�� �� �(�� �� �  �� |�N"�dV�V|�,X�\:�bJ�,D�D,�`Q�6D�0NN���P�<�(��
� ��� �`� `�`� `�`� `�c� `� �0 �
�� �`� `�� �`� `�� �`� `�c� `� �Z�� �� �$� $�� H� �Z�� �� �� � �d�� �d�� � �d�� �d�� � �d�� �d�� � d��0d� �x�� ��	F�� � �d� �2�                                                 �(�(�(� �(  �(�(�()&)Q))  �)�)�)�)�)!*K*  p*              ���0}���������������� ����0}���������������$�����0}�������������������$�0}��������������������
$}�H�$���$�H�$���$�<�$���$�<�$��������`}��$���`��$���T��$����T��$��������T}��$���T��$���H��$���H��$��0}���������������� �0}���������������$��0}����������������$�0}����������������$}�<�$���$�<�$���$�<�$���$�<�$����T}��$����T��$����T��$����T��$����H}��$���H��$���H��$���H��$������  �P�(((�!����                                                                                                                      +  +>+[+x+�+      �����((������m�����������������Z� �����m�����������������H�����$�m�����������������6�����6�m�����������������$�����H�m������������������ �+�+�+,�+� �+  ,  (,M,j,�,�,  �,  �,�,-  :-  O-d-�-�-�-�-�-  �-�-�-�-.N.    �.�.�.�.�.�.�.  m����������������. ��.m�i��m�i��m�i��m����������`m�H�`�HȦ`ȥHȤ`��H�`�H����`m�H�`�Hȡ`ȠHȟ`��H�`�H����`m�H�`�HȜ`țHȚ`��H�`�H�$}������/�������1���m��������������������������������������������� ��`���.���m����������������`�H�`�H����m����������������`�H�`�H���`�$}�����$�����m���������������/ ���m�`�<��H�T��`�<��`�<��`�<���.���`m�H�`�HȬ`ȫHȪ`����`m�H�`�Hȧ`ȦHȥ`����`m�H�`�HȢ`ȡHȠ`�$}������$/�,/ �,/����.M�������������������������������M�������������������������������M�������������������������������m���������������������������� m�`�<��H�T���.`m�H�`�H�`m�H�`�H�`m�H�`�H�$}�����$����� �������������� m�i��m�i��m�i��m�i��m�i� $����� �������������� $����� m������������������������������������������ g/x�x���� [/  w/�/�/�/�/�/    �����((���	����m��������`� �	��m��������`��	��m��������`��	��m��������`��	��m��������`����}��������`h� ��������������
���<1����]�ɛɛɛɛɛɛɛ����P1 ���]��$��Ȕ0���$��Ȑ0�����P1���]��$��Ƞ0���$��Ȝ0����]��$��ț0���$��ȗ0�����t1 ���]�����������������
���t1����]�ɗɗɗɗɗɗɗ���'��  ��(22���]��������0� ���]�����0����]��������0����]�����0����]�����0� ]��������������� ]������ɰɮ�����������ɮɬ����� ]���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          @@H@c@�G�S�S�S�S�ST.TvT�TU!U�U-[-[�`-[�`�h�l�lezez�{|x|�|�~�~}�}�j���N�����������禵�Ѱ�,�,�a�������������                                                                                                                                                 ��p�����	��� �� ��p��p��p���	���
����� ����� ����� ����� �������������� �������2e�����2Ler����������                                                                                  pp  �j�pp ��pp �j�pp ���pp �jpp �jpp �jppp �jppp �jppp �jppp �jppp �j�pp ��pp �n�pp ���pp ���pp ���pp ��pp ��pp ��pp 
��pp ��pp ��pp ��pp ��                                                                                                                                                                                                                                                                                                       j�̪����z������̺z��������j2EeVeUDz"""24EUzVfvUeB3kݼ�����        ��� Ա .�� 1��L?A��L�O�lL@� /�� �Ҳ��A��!�߲��,���I!�L�:]�M� M��>= 0 � �2�����?�NĢM� 2���/��_����"\�� 0�/�L<�����> �0P��Z!J] �1� L>��.�M/�"���-M/��;/� ݲ=!�A�[�� "� ��O��  ��=. ���Ĳ�>/�= �+  �;1����� N����2�����>/.�� �  Բ�C�/���0�<N��M ����0��. .�������/����L�� ����
�� ������ ����/�K������ �#��..���?�/��!��] ��Ѳ�O!�O��>/���
�N.*#���M ղ�.//>�l��<������N/��N �� ����.ղ�}-\��@ �������->"N��1�#����-�M��-��l0�� <�_.1��._���L>;?/��#�B��  .��,>�l�<����Jn���>�N�?��  ��1-�#�.! :��0���.�]��M���]���;^��>�C����O��-��@��}~����q���¢M�L���N^1/�/����-Z�$�B,���r�\��������+0 � ^�-O��@ �� *���<  �>�<^�Nb���!�/,� �/��+\-��� ��-N��@�����#��[�.Q��/�@�����K?Jխ�\"���3����!��!���
1����0������<=> ��/�,^������/��K�-!��/ �  P��,��-O��/��.��[ � �?�� ����<�=��ѢN;5��� %����+Ҳ����/����z��N�����,0����=�"�O��� ���2�Q���C|� �=.�^�����L��_��/O���>� �K[��/�/�c��^.L��/��?���Ĳ��m. �A�@�M.� �l���B��"1���+�! �M� ��/"��0�� > M�"��.��+��"��#�O�;��>���R�>��<��ֲ���$� ������/� �;2���i?��+�"�M���l��{�:P����1� ����?\  �Z�1-2�2�������M0����J��-��!�Yþ?���-�/�N��� ��]�/������ /��������B�1N?:A�����>�[��//m2�[��1�N+1J���� �>�����  ��o���;�2=�����W�².'�`�/���=�L��> ��/�/N�в�/,����Y�}�4������.���< -�.� ž]!���>��1�? .�;  �=2�?)Q޲?�/�0������-�N �!�+.��0��, ����>���>�<���<���+ ���/���!< ��\���-�Ų� �� 1/��  l.B��!�p!�����0��1K���N^���?-/� ��?��� ��,���=AҲ�����*\�#����Q�A� �J>���?������Ol�K�/K?.Բ�-����3�O���\���>������N�+^����������*���Z0?֠�B . ���� Ա .�� 1��L?A         ���L�/  �  o�P �[����δ�= ��ߴ  �" �  -�?.���D0 ������-�� �L�L¤�  $� �d��0#�C����!��-�    �����Z�O�����1�.���6M�P ���D���1�Q��.�:16@��V$��T�`�������� �"��O����C���� �p���%+Q���  ����@��T� �2���#��!� " ��=�3� ��e;�����.�o��@?�0����_�" �<��Q��c�2�� 2���"��/ ��4��"��ѨQ��R���#5��1��S���.̤��4*�B�C>�/<Ѥ�@���4�#��C�!��0��.ݲ�> ����� ,�#�ϨC�B���R�\R�C��ޱ3/���-�B��>���B���?���D�@�!���O!��#��� � �3�����n��:��G��.�5���#���Rݤ ��N���-�C-���,�6?K �D� ���1�$<��Ϩ 1��3�/�����Τ�.�"2���?� $�� D����$��b�C��� ���-�$ޘ��d��<5���C���2���4��-�-! �2C1�F4Q��p�B/��&0����;��o����O��Qβ 1���"0�R���B�/5#��s��B ��2�CИ��.���A�-�# ��Q��� ����$^�?.����#ވ�E
�U݈�p�A���Rܘ�$��0�� ���T���Q�/��%�� ���"�� ��� ����D߈�1��s���@�A�  ��1���@Ј! ��MΈE�2��"��3"��D.������2������ �$��"�2���E�!�3�3�e��0����"����2$���Q��42���3�$�A���5���4 ���߈#A�� ��xCB�U?����D ��$0���!��� "1��xt��#e���E1��!�/��! ���x�"O�����5Q��D�C ���D2���41�����EN�����  �� �x�t���Ce=tm�B4UBx$1 �"��"������#/���x��4R�"x2��Ed?ۼx�UO���xT��D�� x!���4/x/ͼ�FT���"" �ha�t �� x���xR��DC���  $C"����3"��x3�ܽ�x����$x3�1�"xʭb�h#S��dC2xܰ5B�x��ݼ�FB�0��#1��x"��31��#41���2"x.��� ���hd
� ��vx0��$2��x5D��h��&D��3X=/NO�M*x����h����$#hCc �x3T �4�x�����x�$!����xER��3 h ��15Qx��FQ��xD���h���b�x����x��$D�h3R$#��x�#�����hܮ��x�1 "Cx��"!�x�U@��!x��4 ���x�޾C/�h��3O��5ehb@,��e!h#50���x"����h� �!Ch/"3Rx$���#xC��X���/��x��D���h%D@"hRB 7UAX������x��!1���h����Ah/"!edXD�ffTDhۮE0���X���A��X�`ڜ���X!!\L� Tx �41h�!" ���x������h3�̬�3Rh ��FeTh2 ��V2�x�����x!"���!!h�����4Ch��$vB.�h� D"hA���h��������X�����"3h32�Wdh"%4!� @h0 �ݼ�� h������X�3��2B=h��3 hC02!!h4��2h�������h���!��h$C"!1h""$#�X�͛��h������h�TB0X�Fco�RX��$ue%h���2 ��h�������X��ï��4ch�"#D"h22 �h����X�>��Ϳ�h� �X412&C�X��AP �X�#.�0X�ͼ���X��ښ��fh2�$" h#D� C2X�̜���h�������X� "#h!43��X2Q2���H#c����X������X������h�$3!!XQ2"C3 X����>Mh����X���$cSh�4S2"�X�gd?̾�h���X�� ���Xݿ� `=��X202EC1XAeU$#��X!#ξ���h�����X�$�2` h�$X""��X��ݼ��X!.ٻ�##X �����1XBQ4��XV3  "2 X����ﭭ�X����X2�� 31X CE5#H2aEP A�X������X������X�����&DX��#3"BH@1BAUduX�����X������H��3UB H24g#�UUH��!?!�H��̚����X�����H0!C3H��&��HEC���H�������H��������H�� 2S0H32AB@  !8CC ,� !H ���� �8������8��D4"��8CUB���(>RE%/�(��.�(ޝ���(����#PR(2C"B#"!("C1 ������ΐ����� �����#T@  @ #�     ���        �����#4DD�L�ffgvff�333323�ܖ!������������#4DD�L�fwffgv        ���������N jD "4DEfg� ?^���������N         ��7zC"#"#33DzEUfUfeDTzC2#2"33DzUTfeeeTDzD"3"#3#EzEUVfVUUCzC32"#334zUUfUfUUD{332"233D        z�b"#"!J�������3� ""#!0]ʴ/� � �%�   z!!"23DU�"4C42@^ʴ/ �   �	�������j�������#�  �=j�12!���̊%� JС�����3� ""#!0]˴/� �         � �    � fʡ4DEg�   "̪�fv��#4E���#Eg�jO""43ED� ����/���  �    �z�]  !�333EU��݊_�  �"""""�"z"13#34D4�  ������������      �          �?"����/�@ ���=�/�����@�pU�հ� �N�2�"���.�@��P�#��հ�@�P�S߰��=�A��!2����0�!��1�����>�!�0�#���,��O�0�N�"��2������=� �-��a�"�[�5��"�\�� �M��1N���1>���0�>�� ��<��A�K��5�1�;�4��2�+ 2�1�� R���"`ӾM�ү=!� �2+Ѱ%��!B�¬LѰ�1�*�$����n#���0��%�н2~1����/�:�B��"\�1��� ��+!P� ñ3�<1-����
_ ò�?J�%��	!mᰢ�0J2����1[!���/�K �@��Ġ"; ������!]Ӳ��?�J!� ���,0)#�� ¡2K?�:%� ��!�KA*�� �ү!K@*��ѡ"<@�;"!���ð?<1>����%���!L  �$�����2+?� �����?��2M���#����#�L��ck�	��"� �3�?�-!?�� ���/��2=�0�1�������2M�!"����/�- ?�$��'�/Ұ�2< #����#-/�+! �����N�IQk����A�z ��� ���2z0<Ӱ����<�����</�Ҡ�� j ����+?k��ғ�� ��, >����L ����I>;\����M/�L����J�.> ������,i-Q����L.;�����+/n/����M�2���M�>����=�a���J�.������[A�����\ =���=C��� o?���.� ����,@���^ ?����.�5��>�1���P� ^��+ -����W�$�JQ��-�p�O���<-��������D��>�Q���O�����^�?p��a�_�p�P�N�,���=�.p����>��p--�lp�M���?�=p��,!�p�n�=���=p>��O�?t��
!�p�@�/��=`�o��`�0p��N�0�`�O�0��`�@��P� `�.�P�2�-`�A�>�0`��>�P� `�.�B�"� `�3�� �P��/�PO�$�P�M/��PA�1�! @�@�e�#�@��?�-�@%..��O0�1�m�Q�#0�"���.�0��<�>�-� _��!� ,��L�O�\�r���$ @�� �                       ��/�3$����! �1����T� �Ƣ!��#=��-�3��2����N̿�@� �C��� ���� !�����/�=�#��4���M��!�M��%��3��q�$���bB��3��W��0����oT��]�c��k�M������C�TN�S/Cʼ����"��"#��"���/$2�m"�� -��!0��!����.M����C54� ����� Cf�B�������@ ����� ���2��QC��U���+��� #��2 �!�� �@� C2�Aۦ����^�c�> #���P��/�""�+���IU���ND�.N� ��ж�� K3O��2����=�3 <3P��R��0�$�"-A�c�!��0$��M�Q�DP������@J��1L����,.��1�P�S�� ̯,�_�!��P�$�����P��B�?۶���Q���P��O������r���@��b��!�⽶E���_�3��/�����1��n�R���?������" �O�A� ��O�����$���0�C�1��P������ �D��1�����@�� �4� ����P� ��R�C�=�N���2^� �3~���н3]�2�Y���J_ⶬN>�R��3��0ᤶ�O >� 2.�#�� ��@�1-F����./���;��.T<��� ��.��2�SO��������m��a �b/ܠ���0�1�"0�a +���� �!�0�B�b�K��ݶ")��O2A��c�\���� �.#P�%�N�����1��o ��>����Q��#�,/�����!��� �����!����=��=����#����]�e�,�����#��/�����@�� ��Ъ�_�-����2!���=0�޺P����O=�� ��B��.!�� �.�4�aO�����/3��A�@���<�  $�!1�� ��/ � $/� "��J��"�"��O!���<����.�2��!����L�0���J=�����d���0���>�O�S���!"����0�!���$�=�3�����4��� �?�#��2��N��1�A�����N�S��B�3��/���.�A�C���� ���A�D��@����/�S�#� �̲"�?��?�e�#κ�,>���5�.���@�#�  �� /��/�  �//��",��M �@�001-��-1��_�M��϶��A�.�02N�� ��1�� !.�����
$A���-���]��&0����0 �� O����?��� ��O��/�@Ҷ �!�� /ܶ.�o�!�� ��@�!��>�n���0���A�@޶#@�o��0���B�?�3��L�/�/�2�?�32��b@���=��!�.�2 �2s�����>�6.�@�D���� �@�/�>/2������#���2 $�����$���VP5����.��<� @!���@���~�?�K  �=���@�L��-1��2,� ��B����1=�0�Q�0���B��?J�O�\
�Q��a.�ѶP�#�c;�"E;���ʻ�b�T[���#?�������T\��3����$.��3^��3,��/��1��31��3����N$d찶D��#�ݺ,�2���b� ��!�������f���<����#�����/�^���4޶%��`�b����5��?�R�D���$�N�2�B*Ҷ�_��@\� ����@�O_�!����C��@B�����/�$.��C���Ӻ�!��-!>��.���p��$>�/�Tߺ.�>�%O��E� ����#��A� 6������,�B���FCC4����.�D޲�WTe3����E��������"�E����%M �����@��A�"�O ������2�.�0 ��� ��2�/�� �,�.�!��?� �0��N�/�2��O��1��@�0�1���.�C�B��!�"��?�C�Cܶ ��/���?�S�2����A�n��0�E�"�ު�=J[�-\��%�/��϶@�#�  �� /�?�  �//��",��M�?�001-��-1��_�M��!ζ#��A��02N%�� ���2! �� !.�����
41���1����\��&0���0 ���O����@��� ��@���OҶ/� ��0/ܶ.�o�!�� ��@�!��>�n���0���A�@޶#@�o��0���B�?�3��L�/�/�2�?�32��b@���=��!�.�2 �2s�����>�6.�@�D���� �@�/�>/2������#���2 $�����$���VP5����.��<� @!���@���~�?�K  �=���@�L��-1��2,� ��B����1=�0�Q�0���B��?J�O�\
�Q��a.�ѶP�#�c;�"E;���ʻ�b�T[���#?�������T\��3����$.��3^��3,��/��1��31��3����N$d찶D��#�ݺ,�2���b� ��!�������f���<����#�����/�^���4޶%��`�b����5��?�R�D���$�N�2�B*Ҷ�_��@\� ����@�O_�!����C��@B�����/�$.��C���Ӻ�!��-!>��.���p��$>�/�Tߺ.�>�%O��E� ����#��A� 6������,�B���FCC4����.�D޲�WTe3����E��������"�E����%M �����@��A�"�O ������2�.�0 ��� ��2�/�� �,�.�!��?� �0��N�/�2��O��1��@�0�1���.�C�B��!�"��?�C�Cܶ ��/���?�S�2����A�n��0�E�"�ު�=J[�-\��%�/��϶@�#�  �� /�?�  �//��",��M�?�001-��-1��_�M��!�        :�4#�� J��!1�ZO� !�J�&���Z���T"��Z�1 !Z #1#<j���4e!�j��2" ��Z3�?�"z����%d�j��D!!�j4�%A��� 5R��j��BV0�z���ފ���W@��j�b$A� j3U!뻊 �%A��v?��#4D2j"�܊��� a��� j1$B"!��  �r����  Z���������A����!�j� EVD/��   �B�ݽ�  j������ � ���$�B��� z@� 3""� �����C��� ��� ��� ����듪T�� zA� �3U����۠�F.�� z�����"3���� "���A��  �5B!��$z2ܽ��۪�4/�� jVk�����B��2��GO��vFUT!��z4 �� �ʪ�4/�� z5-�����!���C/˚�F?��!jQ$ ��$Vz4 ����ʪ�4/�� zU-���� ����3/��GN��v�eC"��%z3!�� �ʪ�4/��j������4���� ���V>��jVA� �fz40����ɪ�4/�� j�& ���Dz"˩�۽��WN���!v�4D2��6z30����ʪ�3/��z����"�������4/�� zQR�  4zD �� �ʪ�$ ��zr� ���"�������4/��z�  4zD!�� �ʪ�4��zA`��$������ͪ�5 ��� v�!����&z31���ڪ�3/��z%�� �"�����˪�#0��� j�R"�%gzC0����ʪ�4/�� zB� �"�����˪�#0��� j�b gzD ����ʪ�4/��jr ��E�����˪�$0��  vb��̻�zD ���˫�4��          � n �_�D�ln��� ����n��_��������@1/�ϳ�#�/���-A�N  ���2��#�����<����"$!�������SC4�����0O�ѿ��$$.�������P4��O����ѯ�� ������0� ���������?����N�-���>�0 �C4����<߸[�=��L,�N� ������+P��"���.  -��M��'ew�aP�o��{<�ϴ�`>^��?�������L��?�:���@�N��2@�� �0�-�������@B3�� �"������"��0����0���cC ����C4���/������1$^�����/!22��,���b�!�< ��"R4S4>�������"B5�<�����C�Ҵ�� ��/������,���?<_�!� 1 ��$22� ��@����1?1/���� ����2�����O��������/!�����ݽ���"��O��������2�P�!�A1M������0 ��#�������0���?��/��"�QA�"�����
� u!������� ��2 A �1������/A���&�*1$_�����%&����#%@�
*��0���D/������1! ����#�QC��������!/$%2@, ���/����$3<B����J���C2�����1 ��.���:, �@R������>�!"�\_�/.����=/N�%=����� �/<>?�-����� !_-2���,� ���@�0C ����/��$�1����!%�!� ��<!`�����,�3.�1/�����MN_@��?�-M���#!0J2�/�����A"�����!.#= �>!?@!����-��. ^��>>��.?A�������2�"��;�� !�; ���??nA.�c�C�����M9$���o >�������� �� ,1���A>M ������`�]]>__��.
) N4�����!�3���@�T ��� ��;����?�������/ ���0� ��1_��>�P�]����� >/�-��/�N�����..�����>�� �=�����O� ����L�>�,P_�A���?L�?��/�0�A ���!����2��N0����������� ���>���>_0��*��_��= ����."�,����<�޴O kM$�?�� � �����0@����� #��M�1�������F��N?����! �=[;������ �/����!ⰭJ�@��n� ����M0.�L1 ��?���?�M���1���������?�� ����  �� A��а� /�C�M0��K=�,��� @�I ������*B��Ӱ��2,d� ��� ����������/��4N<��Ű�;: ��_�3$�Zݾ�2oC������0$����������������" 1�,��  �?@�?� ��N!n00�����>#R�������B� ������,$��P4/���M1+���1�"�2 ��@1b����+��������"���"���0ǐ��0\Ұ�@�-��0��.?4>��  .5�0�ݡbn�!��B�� �./M/��  �����0����B� �������>#� ��.���@?ů�	/ �3�ఱ����%�����!�?�OP�?Z�;]�;�^M��]0��?���������#��������� ����� ����>��. ���o�M���� �^C�?��� ?��-���?3�!�� ���?�� �/Q���������/ "0���"O�����3?<��-O��<��:B�22 ���,� �n�+Q!/]հ�O��,� ���]$�>@а /ѽ��3".B� ��O�����������
"Ѱ0�.����-��� ��;A�@�=/�
. �N@+n��Y/�?�0<#���@��! ��
��u����A���������M�!�K�O��-? ��-��=�!/O ����1��ô��[0�ħ��K/���1�����O��c���� !��\���K����!а ������ ����β�!�����=���]��Q�K2@� /����0������3��� �Q� ����"02����,O���A�/�����Z@���!�1�O>.����?@��_���������?/� ���/�� /�4Ds��[�۠ ���_M1�  �<�/���ZT ?�/�-3����1!/�0��� ���3 R .�����!���!=B�"�?��/�E۠��� !�_0�?�Л�1���E !>�����2��! !�02��ߐ�/��!�/�- ��! ���;��R�]A&�KА-[�0��^!/;��@�AQ�+����,#�=1��,��� .�3Ô�����>�,��" ��B������2��3B��ۯ��O3�?/������>"!!2��<����>��.. �A.��� �� 02P�+^��/���M� M6�O����-�@/? �=5������C^��O�C�9� �.1���O �L���>B � ��p�c� "�����Ap£��m1 p���N�?c$p �*�?$�p!>>�?p���#Cp2R-�?p�����N!p���.�p�* �pPP� ��`��2$B�` � �/�`���10` ���._0`��.."` �//��`��?�2P>�	���P^���� P�����.bP�Ҳ��!@��<���P  ��>�@��L��#Q@"����@.=�]!@������4{Z�+  0#�M��$.� ,0-�K��0N#�  >              V       !���r$� ���A� ���A�0����A �/�� �B�0� ��A �0� �B�0���B �!�� �B� ����Q �!����1�1�� �B �!�� �B �!����B�!����B �"���B �!���B �!���B �!���B �!�� �3�a���t/�!�� �B �!�� �B �"���B �D����f�R����e/�C�� �g�C���f/�S۱�V/�S����V/�S����V/�S�� �f/�Dܰ �f/�Dܰ��U �D����f/�C���F �3���G/�C� �f�Dܰ��V?�"�� �$�D����6 �2���%0�2���%0�2���%0        z��5U3 ܊������z��5Vd2z44!���j5VD ����z��ڪ���zET1  4fzdܻ�5ezC/������z̫��#2"z33C41 �z��DUR���� ���z��4Ve2z4C!���jVUS ����z��̹���#zUS1�%fzT��EUzS������z˺��"22z!#444"�{��5UC�        z ���Ff�z�� 
%�.����#1���2!D4?��!!���� /����/B��� �"̊���� ���133/z�$A�3��z������z�33 Fa�z�3/%N��z�ݼ�� �z S1�z$1�S��z��� "��z�41�z" �#3���z������j&UD4zC��4 �� j����0ܼ�z�D! 5zO�C��j����ˮz ��33z�4R jܬ�����z�"B # z��4 ���z��� ����z��C2"3j�e/��z�� ����j�6u2EQ�z�#2  �z� ���j�gc4c�z�3 ��j������j�g$E2�z2�  ��Z�Q�����j�FTEd0��z# ���Z� ���ͺ�jDDVC�z"����j��� ���j%D4VC��{"!���         ��K="� �;]-!������ �������.>�*m�=�N/,0��? �K�A�zn����+ � ??� �0�,�2�_2.���� ��� ������������$d�����iLMҰ��������2z����6�����NQ� ���Ĕ��:��>� B#!#�������N����<.� �� ������ � ���������ɛ��-�,�F1 FU��1#���ѐ����-$�.?��-����/��A2#t��0��]�� �����D�/#��߄���.P�O������`_0�������/0�OB^p �������`�E�o�$�"�α?�4�"��K�P��-#Z~�#����z�P1�td�:/�j�j@@x��>�.�S��_�>9�B�  ��D�� "./�A=���2-�n?K�O���KQ���]0�=-�� �/-$!��3��#�����4��C�$=����,��S�#C��� MBx�0b:<�a^��������  ��^�x������x �@ncф����O����>O[`t���0��tK����t�.C�� �d���4�{d/��$o�h��T��{:tT��4�τ3���x�&�U;�?x�#�$.�0�xT��0�!�"t@͢��Sd"���qt-� � �t�N�A"��t���D���d��s� �t�!�B!t.����@  p� >N�t��*o5��-po�����1��?���=���S��A"���\��2�3�U����#t �2C�K��t<��NP��x���P+��%���!������Ԁ���2! t��?��t>� /��t��01��t��! ���t 2Ӥ�������"�2������� ��N�.�CS�Ϯ��"�Є2<���O��NS9-��[��N�����qa���$���՘N,>��� ΢�$!��!� �B� ��@�}�3��."�"[�"�ј� � ��-�/4��!��v����"<������㤱���&$!�����.O�����#��!�� ���\���<�.�O��!_������"B>����n�������/�1������!�\,�"��B��� �/�� �4!�૴F�����m�?2�=�R���6;�Ͱ ?�B�"��"/��.�B��_���� �C�� ��N  �� 0��0/�3]���/�<�.���A��������� ��4�//� 1��� �� �#3��P�.���>�%O�Q��.%�O,޿#���2��$A��>,�s�'<���"���S1�]␳��LM#����������&����2�.o3�����C1��L����/�L �����@���0"����/�b1����`?����.�!��O>!����C��Cm���4=��V0��"5��B��1 ��@��� � ��1���C���=������1��>��� /��R��C0�������4����3��2�Q� �?���#3�����1  3��"���2���3�� ?��0�;�NP��tG%���"����3��x�=< ��xK#<�?�,t ��!�/p#
ڽ�#Pt �� C.��t��4�3�d����t�62��R�p@���5��������/��/����B�� pܬ�C�5_u��c��T�        ��R���?�#z.�"��z�3��0�O�   vd�$A�� ����L�_��! ���A�1������-��!���  !ߚ���T�/��""�z/��O�A���� ���d���3 �z$4+�3���2�ͪ %`�����C�����" ����D��! �C1���z1  �����#?���-�/� �z R���$��A���b!��3z��S���=����v��#�1���!z��u���L���E@����"Ffe��z��eO����$1���c��z��EA�ݼ� �1���%@� � z���� ��5B��ߊga��j/��#0��ߚ� $T���4S� �j-��"T�����e�̊s�   z!��$ �ݚ��E0˽��D  ��z!� 1�͚ ��50�̚�$B��z �ۚ��41�ˊ�Ff/�� v"���$-���$2�Κ�D/�� jR��4��� 3Aۚ�C0�� z$�  �"�����#2���E0��fS "�$-����%t�뚽�50�� f�C33 ������%d.����41�� f�$"F?��������$d���E1��j����B����d����5A�� jb���D>���� T/����6A��j��"��b����� DA���$B��j�2=�C.���� D���6Q��j3��2����D!���5Q�� j�C �E.����4!���5R��j��3���31z����wS-���&Q�� j���T0��� �41 ���&a�� j��!�CBz�� ��WT>���&Q��#j�T1z����VCR���&a��"j<�#�D2z����6c"���b�� z���3z����DDQ���%R�z ��#!z����#ER���%a��# z�� �" z����%CS���&Rڰ# j���D2z���CD��bڿ#!z� �"!z���DB���b�#0z� ��"z���CT���bٰ#!z����"!z���#U���aڿ#!z� �3z��3D��0�� z�-�"z���3D��1��zc��3z��#D��1�� z� ��2 z���#D��1��z<� ��2z���"D��1��zN� �"z�!��"4��0��"z���2z�"��C��1�� z>=��3z����4��1��z2 �2z�"��#��0��z�� �2!z�!��3��0��z����2z�!��#��0��z����3z���2� 0��z ����"!z!��"� 0�� z�� ��2z�"��"� 1�� z���2 z"�� "� 1�� z�  �2z!��� 1��zO����2z!��� 0��#z�����"!z!���� 0��#z���3z�"�� � 0��zA���Bz�2��� 0��zA���3z�"�� � 0��zA� ��2!z�2�� � 0��zA���3{�2��         J��������J�������Z!! !#CZECT22324Z �����Z̼������J�4dDeEDJa4B! ��J����ʜ��Z�� "4CZ4ET4C2A!J �/�����Z������� J�RS!$Z  �����J��ʾBDSZ�4C3Z&2 �/J�������J������J"1!:mέ�J���˛���Z���4DZC#4"2C2J`���ΫJ����� � J� 2A&#"JCB2O"!�Z�������Z������4Ej #C" J�UD#S�Z������J� >4MZ!20 Z�������Z����1%j5EU1" #Z2" ʼ��j��������Z �"45UZD4FR�# Z����۹�z�����5zT""j�������j˼���� 3Z3CT"$EDgZDe#U"!��Z��ٞܬ��z� � ��#V�D!�  j0������j��˽�� Z2"UFUDDZ1 �D1�Z������Z�!R3!1�$1 ��  Z^���˫��Z�̻ۭ�#j!�!$0Z4���J�D� ��!j"C"C!�z #UQ��Z�ʾͫ��Z�������Z #@�43Z2� ��Z���� $Z!UEgEgTjUTR�Z����ܫ��Z�������Z�� DEU1J@��2�Z�������j"##333j1!"43T/�Z���ˬ���j�����z����#C!Z�#�F!Z͹����j�!34D4TZDDgTCf=�j�������j������ފ ��#E-�����jU������j#D2ETeCZDS$32 j��������j������   ���$�R���@�j�0����z5 $12 Ze#!/��j��������Z����B#"z  ���͊�#A��0�jp�1?��z6RB  ZB!!����j�۬�����Z�$U"5CZ  �˪z����D!!�z�#�2!z$C4@� j�!����j�������Z�"UD21Z!  �z����4?�z��/#"4z""T j�0����j�ܾ����Z�2#e2�j����݊��� 2�zo� �0Qj6cEA "jE� � ��j������  Z�A4t Z/ �ݹ�����E0�z�Q�S�D#jcdB "j" �����j�������Z� vcAZ�0��������!!"�z�f�423z3#2 �z ����j�������Z>""4STc�Z��!��쫊���4>�z��NB3EzBC�"jA�����jݼ��� Z"33CC4#2Z� ���콊����� Bz��0�C$T"z4B ��j%
�̙���j�����"Zt35d !!Z���ۼz������$zd�4"433j2$S���z/�������j����"3ZTVB32 �Z!�����˫z�������6ze!#$T #jBE22���z� �����Z����$CUj2C!" �Z�!����z�������4zUE?�EPBj4"3"���j�����̫�Zݫ�#$CTZDFfA0��Z��̫�z������#zUt�t�"3j3@����j����ީ��j���!#2ZDET12�Z �����z�������5zfCC "j!%2��ۻj����ɫͻZ �"fDUZGc3Z����̻z�������6zeS $B"k %2����         t�˼����߸ 2 �2"xD#33"3!,��/���>�������������>c�,�E?��a�+OA ��/��0���� 0���%3�B��34C33#3x44$343#2� ��B���u����������� �#���"� �@��~������������#ܘT?� 3�ƤS�#1��A �  �2S���4��    �$��  ��5�������x�ۼ�����x�������݈�������k���0��/�U���$/��3 ���0"��!��0� �bܘ%�������x��������h�������̨ >��A���e��TD���!.�"���2o��B�#K�F��A4�x3T4D33D"��]�!Sͨ�0$���T�R�
�-��b��0�"���A�?��!�����"��,�/�0��2��4!��B�Q� �AѨM�"��1"""!�""""�_��O����$���?���Ӥ�"���� ���/� ��Q�"�T���^�U�C��#��"F1�! �$0���]�  !��  �@��� �2D�� �B�� ��� �A��"���F����2�}�� � ��R��"�ߨB����>�0��Q�2��2��-� �0����`��E���Q�"� �U��� ��#���R��!��!��?��A�� ߤ�   $�\��/%@?��5� �/�B���,�]���$-�a  �! ���/�M�3�����/����-�U�� �" ���P���"�3����m�5�!��@� �^�?�=�o�1��B��>�"!�B��5���@��4�2� "���@�¨!�"�#/�����D ���!�5������� �=��,� ��"���@�3�c�
��4�#A�! �P���%<��S��,�R�"�4� �3��$�$�>��3� �� ���O��0��?��>��7o��%����E���"@��!���e��D�o���_�ФU�A����>��$�ɲR�ڠ���O� �B�C�>���<����G/� ��D��/!��.�.��1���C��$���/�"]�1�"��.��A���2�$��f�P޼� �$��� !���!7P����b��g �����$��?�� �����$�3���$0�2���n���U��4���1��C���6�E�3��������Q���"�  �ڵm�2!�����1���d��@�$�0��*��T�!��3�E�P��� �"�#   OИ�>��>�Ř^��/��R��]�� #;���1�1͘s�>�#��O�D��d�^���6O#!�����! �˱�A� # ����>��?�0?���#A���N�3! �"�4�uT� ��b!����/�0��_����C��� �-�U������D�/�C��A���#��S���@�E�B��Q��0�� ��P����4�" /��2��1_��B���.��F��5��C�!�42�!�.�2��4#�$��b��0�@� ���4�И��S����" �_�_�R�0�g� #$>��/�AU�=�4��P�^���$5�3��/�2��#��E�-���A	�T���"� "�#�1 ����D���1��#�/��A��>���A�! ����$,�1��>�+�%=�1�3���4� ��>��#>�K�A��3+��4����?��  �3�#����A��1��3 ����T�#�.�b��Q�ŀ �"�#���T���1@�5�O� /��/R��O�1��t��k�A�>��#� �S��+�/� �˙�4���\���63��#R�e�5�?��~��$>��-�"?��.��"��/�<�"�A����D��� ,�����R ����� ��@�?�o�^��2��� %�3�-���A��51�F�#�B���Q����/�R�x+��Z�� �t�S�1�A� #�"�>���-�A���@�!�x<��S��&����D��a�a��b̈1�S���P���? �/�^���0�t�2�GeA��N�/�=�3�!��� ��2��2��B.��1�L� �-��1?x��0�N���`�3�F�҄?�/%/�at�P4? $�t%S�*�0�tB�/������O��!���E�� �?��<x��=�q҄4 ��]�!x��/�%/���U<�/��#�C��1p3������^�>�,�-�f�0�t�7
�\�T�x0�e��K��@�]��5�t���G���2�4��� �� �.�;�1��� � ��1�� �@�O��A��xA�`�%�x#�O�>���1�4��3� �A���?�."�t�2��0ڈ�@�,��?t���4?�x��,�_���x.�,�'_x�"C��31�t"&^�@��t#�CA�n��>�2�2Є�Q��t�5_��t��m�>��A�$ ��1�x? ��3�Ux��-�=�Qt,��$T���x=�-�`����1�����B��?� t�^�3��&tU=�f��qx�.�!.�B�x�0�3.͈?�  �.t�N�.�"#x�C�Q߽R���B��3� t�$��2!t�1�"��`t��3=�4x��A�!�5.x�� B� �xQ��"-�>҄!� ��x�o�"x;�-�4�t�V^�  ��t�D��R-t�%B�6_t��0>�Bx�C�u�d�Cb��^��t �e�x�/�?�4x��-�@�"t�U����x��!�x�O�#�A�tD0�%$�t� �A�t��/�@!t��"?��0t���$A���tB�� �xP���$�h@���t/�@�!�x��!� t�1�1p=�" �Uh.�� �M�t1� �D��t�O��!��3x��. �!t".�$�5�hI�4/�c�yB�3�$        j���##�az�2��j��B�4R�j���?�2z��D�j����z2�D?��z�����$z�41�� j��1�D�z�#B���j۰U-��z$3S��  �z�!4ܼzET��zU���3zU>���j#u����fz2��zT���Cz��� ��tz���  #z���ez�� �5�z��s�z��5O��z�"�Q�z �$3��zA �z�%/��z $!���z�1���z4$?���z "�� #z�&A���z2��1�z�'b�� zD���B��ze1���6z-���A��zUA��� 5>z���A��EzQ���/O�z�0��ERz��� 1��z� ��4DT�z�3 �zٮ%UD�z��R � ���3"��z�D"�?�z��eC3�̾zE#�?��z�eUA�ͽ%z�0�ɠzUUA��@z�0�1�ٟ3zWb���A����� %za ���B�2����Az���2�#�����Bz���2# ����Bz���#!�z���U""���  �z�0�"D�!���#0���� "���?��51����! "���@���%S��#�/���R݊�U.��0�� ���R�ߊ$F@���A���#�"�UQ���B����-�2%�c���4������#4T���1������"3C/���1���� C#0���2�! 늬"3""���"�z�DgR4?�ފ�!�#1��z5UT3A���1���zD4DS����B���!zVU���!�B�� �#C����B�����D!���T���"���U�B���C�����5d���!3/܊���5U/���#�ϊ�UB���41��� � ��EC���#C��� ����$31�ЊE.������2"���E@����!��$�R�������S���1���1�U/���! ��#���4B���" ��# �����$C͊!��"����e/��!��3  ���EA��2� ��#!� ���ER����1����d ��!����S��݊�FA��"݊�4/��"�ϊ5C��ΊA�� ��D!����C��#�#�2�"�4�.�� �2z!��0��Q���" �z �!�Sڊ��!� !z�/�z��e!��/z��C!��z�6c��2z��F@���z�uB��1���B���ߊ%1�����C �� ��C ��"��$1�� ��$�2���" ��C���C���1�3z/����UAz��VQ��Bz�����TCz��5d.�!���#�z�fA����2��zT!��C���3 �zE12�$C��2���2z $3��T1���C��#!z#1ڽR��#ܽ�Cz��4 �!���51�jE��$#ED���Sz��C"���42 �z� �FB�ܽ�$3݊�# ����U1�� "! �ۊ�4S/�� �! 3��͊�$UA����C1����DT�� ��5Cʬ��5T0�� ��U0۫��#�5C���ER���4�T-�� �%�T����3D�A���T�0���"4S����DC������3E���   5R�����5@݊�  #S/ڊ��C�E1ڜz� #V>�� $S���z"30�"� �#4>���zB1��C�D0˻�!zB ��f��D2���z#��&r��#3-������C  �4/ۼ�!����4! �3�1���"���4A�1����"��S�2���� 0�݊U!�#튼���2��e2 �0�܊��#��F�C1�"ܾ� �0��t�"�"����!���B"�������3��fS ����� ���6e0�������%e2�1��� ���Vb����  ����TT�/������4T ������#T��z��C��#F�31 ��z�V-��'dG� �"��ފ$.��23����A���T" ����A�ܽD2�����CꊾEB�������B뼊CC�  � ��2���3C �  �����4�C  �� ���43j�����.z$̚VS z/��� &����2"zA���E<���3/����� 3-�z�Ue>�3����4-�ъE"�/݊��D��D�2���͊�#C��EC��� ��T��4C������T��S�����S���D���� ��Sz�v/��z���d�z %1��z��R�"z1"!��z�.�T0z�C1�ݪ�z�&u!�z�T"���C���$C ���3��� ���%d ��4� !���@̊�%e@��A�����P�ϊ%fP���S����Bپ5�vQ���4 ����!ٿ4f�b���%0�����5Uc���$1������$ES����C�������DS ����B� "늬�4B"݊�"�1�z�DVTF>�ފ �2��ze33Ebھ� B��#zBEe���T��"!� D����S���3��D0���!�T���"��UA���!C���"��E�S��3��� ��5d���"2����$U@��� #2�ϊ��FR����3B���� ��ES-���C�����$31�ϊD.�����31���5@���� "/��$�R�� ����D���!���" �E/���1��#�����D2���3 ��2!�� ��%R͊!���2���T/��1��#!��E1��1���1 � ���6R�#/���! ����T ��0����C����EB��"��C/��Ί5C.��ފA��!��S!��!���C� �#�B���4���0�2z0��0��`���" �z�!�!C����"�        j   �l/0j�õ���;>j�M.��Z�	-.+33j����N�v��C3D$z����/??jKA�����j�"?O�z+ �Ӵ%z��=;_�z����  z/-��jD/�Ҽ��/jo%_�j���o<sz0���/�z�!O,��zz����-�<z/"���z 1�>`�0����� ""0���zB:�@C4�1�����""$@ܪ�z&4��3BW�0���3/���!���zTf-��3eU���!���"����5��"3�!��"D/���  ����!D ��B#� ۚ�2D/���#23/ۚ��"T/��#2� ۩�3E��"2#/ۙ��2E/��#1�/ۙ�CE.��31#.˚ъ2U.��30"�.ښ�CE��3!#.ɛ�3U��#1�-˪�2V��"2#˪ҊCE��21�.���3V��21#˚�BU��2!�˚�2V���31˚�BV��#0����CU��30ʛ�CE��#0�-���CF�         t�=��SD�x!0��ܔ���Q �B%�}�<�� ��"_9�5���J"�L#��:3]��p�  ��N��e2O�����/�������N�B�%< =�� �N�`�M,�&�@O��N�/��� ��� � ��"���%����� �$-�$0�R��0�/l��5e/0N���������� &��� ������@�/� �����P��B�^;Ք��ұb�ո�  <��$:�:��� 0�1���������1-� ��J_$�:�#���̨��+-A<�.M@��O ���1?�����j�������5O�TD_,������Կ݈,��-����?,�>cC&4�2�09:�L���t�����+���������L?�.M]�1 �22!�B�P. t�>����dհ���
,�d�1l@#"@x� ]��t� ��h�"���/h�N��Ds�,?43@R(տ/c� �"����        z�4,�Q�z�"�B�z�� ������� ��E0��0� ��S���4z" 4��Q�C!��3�Њ ��B!��� ���뭊���1��zUWu�#1�42/�0.�!!�E��Ezr�$A�EC����f����� �����2��Ί5B��5�D!�2��3/���z7A��UV2C���D �����묊�����2&A��""�FR�%1ߊE1��3�/��5T��� $R����! ��ފ��" ���ފDB��&�c�3��!��!�� �!���%R�����501������̊��"��� D0��#Bz�ge���"! �C���!�5A����� $S������ ���" ���̊C0� "zDBFd�D!��U,��D�����4C�z�ʐWv!3��� ��ܚ  ���z1�TS��31��EB�"ފS/������"#"��� 4C���!������"���z�3�@��T!3���"2��C����32���B.��!�뼊� �۬�z�e��!$T ���5R��"!���1#/z�� Df,Ί �!�����#����z�A�۰�$S#0��D�1 �3z���3E3"z���E2# ���4/��̊�#�����z��d!�!�4D1�"z%@�&t"1��� !Cz��2e0܊� "!��ϊ����܊��ߊ5B"!�2z1�26t����Cz-��3 T���22�̊������Ί���" ���zVTE@�#2"� ��3!! ���"!!���/D0�z�dQ��z���!ګ�Ɋ��1���zFe0B $Uz!��1vS1z���ECC���C ���4B��������ۊ��"���z2$e�Fd.��1��3#A z/��5Bdz�3B@�z�342".�ފ�� �ˊ��2 ����z6c2F!&�!�"#Tz���g0 z��f���D������ �����"���z0"e!���u/�z2��U!5?z��R3�z�d#A������! �����3����z2��$1DzB�UEe!z����fR�z��Dc��z 6b ܊��� ��  �������C!�  ��C2���$1  z1��4DS��zS"342�� ��"�݊�� ����z��44U�!��!T1z-��!DAz��%e1��z2%T!��� 뼊��������z����Wu����DD!z��3432z���VS ��B�z���%b�̫���� ����z����4C4�!�� 4C"z�� FTz��#2F@�z3�GuD0���!܊��������z٭���%u�!�� #D1z���$T1z�%e/C/� "#C/�z���E.�̊������z������DF�A���"33z_��! Edz�4!T���U!���! �� ����ފ������C����#S!zQ���5Cz D0TC��""#3 �z��$Aڽz�������͊����� �!���3Cz>��""!1z�2Ft���$C!z�"3��z�����ʭz�����U�!���"D0j � 7u��z2#CUAz�5U3ECz�� 2��z���ܻ��z�ۙ���$fz@캽UD2j�5Sc2�  �C ��� "31j��ES�$�z������������� 3z1���e3Ck�5CSB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��:�
�v����������*�����r�pX�Z�	�	
|	n�|�����	pT	n�~��h� ���@��Z��z���>�d��6�0��"�����t����v�����n�� J���R���@��4���N�����>�������������v�D�����*�����v�6�����~�
d
��,��&H���<D��V�J
�FP��d�� L� P,�L�������p����>zD $�
�
��	<8	����N���� ������d�|��\R�B ,�>���b������*������d���������T�*�����L�~�������z�R���R�l���Z�����4�����B�� � 4��	�����Z��0dj�	�����f ����n����	���
t�(����
���	���������T��^�^���:�42�$8���d�rD�v p�*���n~ �v�"��D����
� �	�rv^�ZHp��*�d���&V��� �n *. �  .& � 2 ��@ p�H �F ��8 ��. �� ������������L�D�������`������������ ����� ��8�������^f�������^ ����������<� �H�������`���z�,�:���h�
����������$����� D����� �������v�������`�����`���N�<�&�������~�F������������P�������������0�~��������������n�6����r� ���lh~�F��.Pz� � *����$��|8����D4�x v��x�@�\�<�H�h�X����������2���4�D��������~����b�������h����F���X���0������V�&�����(�:��0���v�\�����n�j�"��������|�������R���Z��������� ������v�l�H���(�F������"���n�������`� ������
����������.�����������"�������0�d������������D���d�� �����&���t������r�`��������� r�~���J dnx��n�f � �x�r���^�� ��:�r����r���D���b���������F������`�p�����\���8��� :	� ���
^V<z���|�^vv��
jn ��� \��������Z�������b��������^���������T�V ��� Xr�:� \2�n���H	6r
�	��
�2�T �~ ��6Drp����
�0�J>N�88z��H��8&�
V�<��F���p�

R
jx
�L\�F��b4��������H�x���2��J���P
N�	h�	�	PL
��
F�v�L~�j�f�\&.h��J���������b���4Z���l�
P��h��� ���0p��
��
���	�Z	��D	��`	���	* 
nf
��
��P&�f��	��
z^
h
��	6�j�4���\��	�D���� ���B��"��@ ����h�@����������0�>������������������& �X>���
�p *,�j�
	�vd��>�(j�.���������������*����Z������R�b��:�����4������|���x�2��T�h�f�r�n�8�j���l���~�f���� �������.��v�������V�������@���f�����������v�0��f���P���\�b����������p�J�:���������(���T���������6�������F�Z����X����p��R�~�b�*����f����6� ������������ ����^�0�����j��:�T��:����f�x���(���*�P���2�B������ ��d��8L�|��D���d��.�� ����n�<���������L�0���������������`�������h������J�>��J�\��F�:�������V�����:���"�V�z���|�����R�8�N������:�0� �6�D�n���������� �N��b���H������ �X��HH�p��db>�V~�������������8���������v�f�F��������\�������t��� ����N��f�0	L�J
�\���r���:��&��h$�>���
*�p	��B	��	��
���
B �������H��	�
Z
N	�
vt�:
�0Rfn`f�0��
�

�*	�
6,J����j���B�F�@�� | ����$��Z\ ��z `�p	 �
�����	l
�
�.
��	����$ \B�J�Bd4 *.T@�V�~���&���,����������$�>2�
����
TT&�
�����
 
8�	h�	��	��	J	:���
�� �B�$�d�	�:�d��	��@�������&\���

��	8n	�6	T��, �	��8���.�T^	�6�Tr�����vR":��$�
�d��fb� ���*��������`�� ��8 �����������n�����x�\�*�j���n�(�������:�z���:�D��������>�.�@�P��V���>���������b����@������������2�����4����������x������.�6������`�d������h�*�� �������L�2�@�����H� ������8���h��������"�@���n� �"�����^�Z�����J�\�������l���D����������@ X���0��� ��x�(����V����V���������h�������Z����\��8�"�<�:�t�~���,���z�����������"��������f�J��������4�����$���&���D���n�������������*�p�b�B����>�����N����"��B�d�\���|����^���$�������4����N�t���v�<���������`�V����Z������R����f�����<�H�����X�������@��r�����~��������$����X�|��Z��������H�\P���,�z"�d�����>�����(��Xj�����r ����������B������������V����j������R �� 
\                    �(        F���:�1�������:���	�j� +Y/�+   +Y/�+v�fІІЖІЦж����������� J�  �(�,�4�C�    G�Tхљѹ����X�xҗҹ������	�;�  YӏӦ�������'�  F�tԙ�������+�  C�nՖկ���%�b�z֮֓֟�����  �  ���-�5�  @�  U�l�p�|ׂ׍ר�  ��������F�tآ�  ����������  ���������`���� �%��?��`����
��`�����v���
�`����������  ��������=����m��=�`m� ������H�m�`��������=����m��=�`m��������=����m��=�`m����}��H�}�{�	|��~�z�x�v�w�x�y�z�{�|�}�~���������K��{�|���~�z�x�v�w�x�y�z�{�|�}�~���������=����m��=�`m�����	��=����m��=�Xm�������ɫɫ�ɩ�ɫ�M��-���� ��
����?�ɦɦ�ɤ�ɦ����������
�`}��$�$m����Ȫ�`}��$�0h������������`��@�y�z�{�|�}�-�ɲ�����{���+���
��0m��$����Ȫ�0���(������-�ɰ�ɮ�ɰ�M��-����ɰɰ�ɮ�ɰ�M��-���� ��
�0}�����0�����������ɫɫ�ɩ�ɫ����������
�`}��$�$m����ȱ�`}��$�0h������������`��@�y�z�{�|�}��$M�-����}�m�}�-���
��0m��$����ȱ�0���(������`��-���������`����������� ���
� }���0� ���0� ���0� ���0������`��-���������`��������������
�� m����M�=�����`]�����������
m�k�h�i�j�k�l�m�3�`��k�h�i�j�k�l�m�3�`�� m����M�=�����X]��
���`� m����M�=�� m����M�=��0m�� ���
�(}��0x�(}��0x�(}��0x�(}��0x�����	@�]�=�����'�`]����
 m����M�=���3�`m����m�k�h�i�j�k�l�m���-�� ]��������m�k�h�i�j�k�l�m���-�� ]������������
m�k�h�i�j�k�l�m�3�`��k�h�i�j�k�l�m�3�`�� m����M�=���3�Xm�����@�]�=�����R�`]��^��s�`m� ������������
���Y��I���i��I�����o����$�M��o����$�M��o����$�M��o����$�M������s�Zm����0������`� ����
����;����^����To�M���
�<m����0��H���X����0������B������� ���
����;���^����To�M������<m����0������`��
�<m����0��H���X��^�$m�-������$m�-������ �����
����Y��I���Y��I������]�9�K���\�9�K�9��]�9�K���\�9�K�9��]�9�K���\�9�K�9�� o�O��o��M��� o�O��o��M��� o�����M�������	�$m�-������$m�-������$m�-���������$m�-������$m�-�����������`m���� �%��?��`������`m������v��`m�Z�`����
�`���� �-�ɫ�ɩ�ɫ�M��-���� ��
��0}�����0����� �����-�ɦ�ɤ�ɦ�M��-���� ɦɦ�ɤ�ɦ�M��-���� ���m���$��ɇ��������=��$�m�ɇ������� 0}�����0����� =���$�m�ɇ������� =���$�m�Ɍ������� `]� m����M�=�� m�k�h�i�j�k�l�m���-�� ]�������� @]�=�����  m����M�=�� m����M�=�� @]�=����� ���$m�-������ `m�$�-������ �
m��������������������������� Y��I���Y��I�� ]�9�K���\�9�K�9�]�9�K���\�9�K�9� ����$m�-������ �
�<m���� �
m������������������������������������ Y��I���Y��I��Y��I���Y��I�� ]�9�K�9��\�9�K�9�]�9�K�9��\�9�K�9�]�9�K�9��\�9�K�9�]�9�K�9��\�9�K�9� To�M��To�M��To�M�� Y��I���Y��I��� ����.�>�N�� ��  ~ܝܬܻ���      ������������    	�%�?�S�x݌�    �ݰ�����        ������&�      Tކ޷����$�    (�R�wߠ߰���    �������        ������  ��((�
���`}�� �
����T}�`��
����H}�`��
���$�<}�`��
���0�0}�`�`}�� �T}�`��H}�`�$�<}�`�0�0}�`��
���<�$}�`�H}��0��H��T��`H��`�`X� �T}�0�$�<��H��H��`�`X��H}�0�Ȗ`��H�`�`X�$�<}�0�<�$�`�$�<�`��	�}����}���0�0}��T��`�0ȝ`�`X�<�$}�0�`Ȝ<�$�`�`X����!��,��!� �7��B��L��B��V��b��m��b��x����������!��,��� �7��B��L��0���H��V��b��m����x����������H}���H���`�H���x�H}���H���`�H���x��0}�$�m�T}��0�$�m�T}��0�$�m�T}��0�$�m�T}� �0}��m�H}��0��m�H}��0��m�H}��0��m�H}�$�0}��$m�<}�$�0��$m�<}�$�0��$m�<}�$�0��$m�<}�������_�]������������������������<���`�<����H��`������0}�$��T��0�$��T��0�$��T��0�$��T� �0}���H��0���H��0���H��0���H�$�0}��$�<�$�0��$�<�$�0��$�<�$�0��$�<�������� ��-�����<���`�<����H��`��������!��,��� �7��B��L��0���H��V��b��m����x������� �0}�$��T� �0�$��T� �0�$��T� �0}���H� �0���H� �0���H� $�0}��$�<� $�0��$�<� $�0��$�<� _�]������� _�]������� _�]������� �0�$��T� $�0��$�<� _�]������� _�]������� _�]������� �������� <}����H�� �� H}���H���`�H���x�H}���H���`�H���x� _�]������� _�]������� V�F�f�� <�  v���������  \�}�������    ��)�D�_�l��  ���
����� �
����� �����	�`��-��������0�`������`��-��������0�`����T}�������`�0�0}��
��}���}���}���}���}���}���}������`�<�$}��
��}���}���}���}���}���}���}���������  �_����
����� �
����� �����	�`��-��������0�`������`��-��������0�`����T�}������`�0�0}��
��}���}���}����}���}���}������
���� �
����������	�`��-��������0�`������`��-��������0�`����T}���,����`�0�0}��
��}���}���}���}���}���}���}������`�<�$}��
��}���}���}���}���}���}���}��� ���� ���� T�� ���� ���� T�� 5�  E����9���K�������((�(��(���=��]�=��]�=���]����H��H�=��]�=��]�=���]�`m���� ����`m��=��m��]���`m��=��m��]���dm�`������"0
���
��=��]�=��]�=���]�HH��=��]�=��]�=���]�H��=��]�=��]�=���]�`m������,
�����=��]�=��]�=���]�HH��=��]�=��]�=���]�H��=��]�=��]�=���]�`m������2�����=��]�=��]�=���]�HH��=��]�=��]�=���]�H��=��]�=��]�=���]�`m���������=��]�=��]�=���]����H��=��]�=��]�=���]�\m�������T�M��` ����=��TM���` �����=��dM�����
y�z�{�|�}�~�P����Z�M��` ����=��T���` M�����=��`�����
w�x�y�z�{�|�}�<�� HH��=��]�=��]�=���]� I��9�	�)�� ��  Y�d�r�x���    ��������#�    B�T�w����    ��������  ��    ��              0}�������� ���0���0��`m����`��}��0���0�`m�����}��������������������
d}��0���}��0�`h� ����(P0}��0]�0}�`�0��`h�����F`}��(�0m�0}�`m�0}��`h�����Z`�0��`�0}��`h�����
<`���0}����`h����P�0}������}��0�Xh�0}��ȯ��ȯ��Ȫ`�� �0}���0���0���0���0���0��`��`m��������0�}������0�������������������ȩ��`m���������}����Ȳ������Ȳ������ȧ��`�X�0}���� ��`��`���}�������������������
d0�  �0}���0�� 0]�}��`m� :�*�Z��  �  j�}������      �I�f���      �����          >�Q�w����      ���]����������� ���m������������������������������������m���ɺ����ɸ����ɺ����ɸ����m���ɵ����ɳ����ɵ����ɳ��m��������������������%��  ������$m���$����H������� ����$m���$����H�����������$m���$����H�����������$m���$����`����m��@����@����i�e�f�g�h��i���j��k���l���m��o���������]����������� ���m�����������������������������������m�����������������������������������]����������� ���m������������������������������������m���ɿ����ɽ����ɿ����ɽ����m���ɺ����ɸ����ɺ����ɸ��m���������������� �������� ������������� -��=�M�]�m�� �  }�����      ����            ��?����      ��B�������    ���%�5�G�X�    f������    �	���� �	���(��	����0�m�����`��	������`��	���8�m�����X���P�(����  ��2((�	����� �	����(��	����m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i��� �	���(�m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���0�m��������`���H���H���`�8�m��������X��	�m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k���i�m�i���k�i���l�i���k�i������ �	�m�i���k�i���l�i���k�i������m�i���k�i�������k�i����%�0�m����6�`����0�`�0�m���0�$��0����0�$��`����0�H���`�8�m����6�`����0�X��	����`�����Hm���`��i�����������������N� i�����������������_�0m��$�`���H�`�`h�m��H�0����`�8m����`���H�X�`h�0�m���`��k������i��l�i���k�i����p� �(�`}����`m�����X}�`���`m���� m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i��� m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i��� 0�$��H��� 0�m���0�$��H��� H���H��� ���������������� m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i��� ���������������� 0�$��0����0�$��H��� ���������������� ���������������� m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i���m�i���k�i���l�i���k�i��� ����� ��  ��
�,�J�        V�    e�        �r�Ȇ����� ��d-����������������������������m�������������������������������r������ ��������� ����  ��(PP���m����� �����Ȇ��� ������������������������ ���������������� �m�����Ȇ��������Ȇ��� �����Ȇ��� Ȇ��������Ȇ��� B��"�2�� �  R�t�  ���      ����������      �����/�Z�      _����������    �
��d�<�� ��0}���#�0���H� �
�d�P��Hm���������
�d�P��
��7��
�d�P����0}���#�0���@�0}���#�H�� Hm�����������H}���������7��0}���#�H�@���b�� Hm�������0���
��0m��0��0��0��0��0��0�ɡ��m�0�ɣ0�ɡ0�ɟ0�ɤ0�ɣ0�ɢ0�ɡ���b������  �<�((��
�����m����
�	������`}�0� �
����m����
�	������`}�(��
����Y�0}��`�0��
����
3�m�
�	������`}�0��
����3�m�
�	������`}�0��
����Y�0}��`�0� 0���0��H�0��0�� �m�0�ɡ0�ɟ0�ɡ0�ɦ0�ɥ0�ɤ0�ɤ0� 0}�����0������0��������H� ������� ��  �����0�]���������$�>�^�~������������A�l��������
�d����������0���H� �x�� }�������������� ��������������x�� �}�������������� ��������������x� ��}������� �������������� �������x� ��}������� �������������� �������
�d��������������
�d���
��m�0�ɡ0�ɟ0�ɡ0�ɟ0�ɟ0�ɟ0�ɡ0��
�d����������0���@�����  �<�((�!�>����������Px�}��� ���0}������<��������������0}������<���$������������0}������<�������������� $�0}������<�������������������Px�}�����������Px$�}������ �����Px*�}���������H�� �� }�������������� ��������������� �}�������������� �������������� ��}������� �������������� ������� ��}������� �������������� ����������������m�0�ɡ0�ɟ0�ɡ0�ɟ0�ɟ0�ɟ0�ɡ0�������H�@� 0m��0}��� 0��H�0��0�� Hm�� �0m��0��� `�� %��5�� �  E�j����������  ?�a�p�����      �����������D�  ���((�P�!���0}���������������� ����0}���������������$�����0}�������������������$�0}��������������������
$}�H�$���$�H�$���$�<�$���$�<�$��������`}��$���`��$���T��$����T��$��������T}��$���T��$���H��$���H��$������((�P�3��N�����0}������ ���0}�����@�����0}�����<����
�0}�����8�����0}�����4�0}���������������� �0}���������������$��0}����������������$�0}����������������$}�<�$���$�<�$���$�<�$���$�<�$����T}��$����T��$����T��$����T��$����H}��$���H��$���H��$���H��$�� ��x�x���� l�  ���������      !�?�\�y���      ��              �	����X}��X��X��`� �	����X}��X��X��`��	����0}���������	����0}�������(��	���
�X}��X��X��X��	����`}�X�P�H�@�8�4�0�`� �	����`}�X�P�H�@�8�4�0�`��	����`}�X�P�H�@�8�4�0�`��`}�X�P�H�@�8�4�0�X��`}�X�P�H�@�8�4�0�X�����((���	�����  ��{��|��}��~�����~�y��z��{��|��}��~��������������������`������M��0m��'��9�Z�`� �M����������0m� Ƚ$�M��0m� �M����������0m� ���~�y��z��{��|��}��~���	���� ���~�y��z��{��|��}��~�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   <�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    a��  ` �
��}  `  !"E��
    +"_
��U    +Z���   � 	���     < ��
��     � ��

��    � ��p�z�R�����f:��Yoj��  ���,������f�X!B���[�� } 2	�j	^���� >�+j��  �8��+6)�6�b�@��J���b[U  U 0�
z�x�������f��<�h�0A�H��  ��������������R�A7�l  �     ��� ���%f;�2�%p;���eD8h  �    ��N���h˰���6����� �D�>�g        ��\ #��8��i�X^����   @�n�
   �    �< �l�z�� �  �  ��(<a���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                